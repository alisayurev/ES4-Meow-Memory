library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;


entity one is 
port(
    clk : in std_logic;
	address : in unsigned (14 downto 0); 
    rgb : out unsigned(5 downto 0)
);
end one;


architecture synth of one is 

signal addressOut : unsigned(14 downto 0); 

begin
    process (clk) is begin
        if rising_edge(clk) then
            case addressOut is
			when "000011001000111" => rgb <= "000000";

when "000011001001000" => rgb <= "000000";

when "000011001001001" => rgb <= "000000";

when "000011001001010" => rgb <= "000000";

when "000011001001011" => rgb <= "000000";

when "000011001001100" => rgb <= "000000";

when "000011001001101" => rgb <= "000000";

when "000011001001110" => rgb <= "000000";

when "000011001001111" => rgb <= "000000";

when "000011001010000" => rgb <= "000000";

when "000011101000111" => rgb <= "000000";

when "000011101001000" => rgb <= "100110";

when "000011101001001" => rgb <= "100110";

when "000011101001010" => rgb <= "100110";

when "000011101001011" => rgb <= "100110";

when "000011101001100" => rgb <= "100110";

when "000011101001101" => rgb <= "100110";

when "000011101001110" => rgb <= "100110";

when "000011101001111" => rgb <= "100110";

when "000011101010000" => rgb <= "000000";

when "000100001000111" => rgb <= "000000";

when "000100001001000" => rgb <= "100110";

when "000100001001001" => rgb <= "100110";

when "000100001001010" => rgb <= "100110";

when "000100001001011" => rgb <= "100110";

when "000100001001100" => rgb <= "100110";

when "000100001001101" => rgb <= "100110";

when "000100001001110" => rgb <= "100110";

when "000100001001111" => rgb <= "100110";

when "000100001010000" => rgb <= "000000";

when "000100101000111" => rgb <= "000000";

when "000100101001000" => rgb <= "100110";

when "000100101001001" => rgb <= "100110";

when "000100101001010" => rgb <= "100110";

when "000100101001011" => rgb <= "100110";

when "000100101001100" => rgb <= "100110";

when "000100101001101" => rgb <= "100110";

when "000100101001110" => rgb <= "100110";

when "000100101001111" => rgb <= "100110";

when "000100101010000" => rgb <= "000000";

when "000101001000111" => rgb <= "000000";

when "000101001001000" => rgb <= "100110";

when "000101001001001" => rgb <= "100110";

when "000101001001010" => rgb <= "100110";

when "000101001001011" => rgb <= "100110";

when "000101001001100" => rgb <= "100110";

when "000101001001101" => rgb <= "100110";

when "000101001001110" => rgb <= "100110";

when "000101001001111" => rgb <= "100110";

when "000101001010000" => rgb <= "000000";

when "000101101000111" => rgb <= "000000";

when "000101101001000" => rgb <= "100110";

when "000101101001001" => rgb <= "100110";

when "000101101001010" => rgb <= "100110";

when "000101101001011" => rgb <= "100110";

when "000101101001100" => rgb <= "100110";

when "000101101001101" => rgb <= "100110";

when "000101101001110" => rgb <= "100110";

when "000101101001111" => rgb <= "100110";

when "000101101010000" => rgb <= "000000";

when "000110001000111" => rgb <= "000000";

when "000110001001000" => rgb <= "100110";

when "000110001001001" => rgb <= "100110";

when "000110001001010" => rgb <= "100110";

when "000110001001011" => rgb <= "100110";

when "000110001001100" => rgb <= "100110";

when "000110001001101" => rgb <= "100110";

when "000110001001110" => rgb <= "100110";

when "000110001001111" => rgb <= "100110";

when "000110001010000" => rgb <= "000000";

when "000110101000111" => rgb <= "000000";

when "000110101001000" => rgb <= "100110";

when "000110101001001" => rgb <= "100110";

when "000110101001010" => rgb <= "100110";

when "000110101001011" => rgb <= "100110";

when "000110101001100" => rgb <= "100110";

when "000110101001101" => rgb <= "100110";

when "000110101001110" => rgb <= "100110";

when "000110101001111" => rgb <= "100110";

when "000110101010000" => rgb <= "000000";

when "000111001000111" => rgb <= "000000";

when "000111001001000" => rgb <= "100110";

when "000111001001001" => rgb <= "100110";

when "000111001001010" => rgb <= "100110";

when "000111001001011" => rgb <= "100110";

when "000111001001100" => rgb <= "100110";

when "000111001001101" => rgb <= "100110";

when "000111001001110" => rgb <= "100110";

when "000111001001111" => rgb <= "100110";

when "000111001010000" => rgb <= "000000";

when "000111101000111" => rgb <= "000000";

when "000111101001000" => rgb <= "100110";

when "000111101001001" => rgb <= "100110";

when "000111101001010" => rgb <= "100110";

when "000111101001011" => rgb <= "100110";

when "000111101001100" => rgb <= "100110";

when "000111101001101" => rgb <= "100110";

when "000111101001110" => rgb <= "100110";

when "000111101001111" => rgb <= "100110";

when "000111101010000" => rgb <= "000000";

when "001000001000111" => rgb <= "000000";

when "001000001001000" => rgb <= "100110";

when "001000001001001" => rgb <= "100110";

when "001000001001010" => rgb <= "100110";

when "001000001001011" => rgb <= "100110";

when "001000001001100" => rgb <= "100110";

when "001000001001101" => rgb <= "100110";

when "001000001001110" => rgb <= "100110";

when "001000001001111" => rgb <= "100110";

when "001000001010000" => rgb <= "000000";

when "001000101000111" => rgb <= "000000";

when "001000101001000" => rgb <= "100110";

when "001000101001001" => rgb <= "100110";

when "001000101001010" => rgb <= "100110";

when "001000101001011" => rgb <= "100110";

when "001000101001100" => rgb <= "100110";

when "001000101001101" => rgb <= "100110";

when "001000101001110" => rgb <= "100110";

when "001000101001111" => rgb <= "100110";

when "001000101010000" => rgb <= "000000";

when "001001001000111" => rgb <= "000000";

when "001001001001000" => rgb <= "100110";

when "001001001001001" => rgb <= "100110";

when "001001001001010" => rgb <= "100110";

when "001001001001011" => rgb <= "100110";

when "001001001001100" => rgb <= "100110";

when "001001001001101" => rgb <= "100110";

when "001001001001110" => rgb <= "100110";

when "001001001001111" => rgb <= "100110";

when "001001001010000" => rgb <= "000000";

when "001001101000111" => rgb <= "000000";

when "001001101001000" => rgb <= "100110";

when "001001101001001" => rgb <= "100110";

when "001001101001010" => rgb <= "100110";

when "001001101001011" => rgb <= "100110";

when "001001101001100" => rgb <= "100110";

when "001001101001101" => rgb <= "100110";

when "001001101001110" => rgb <= "100110";

when "001001101001111" => rgb <= "100110";

when "001001101010000" => rgb <= "000000";

when "001010001000111" => rgb <= "000000";

when "001010001001000" => rgb <= "100110";

when "001010001001001" => rgb <= "100110";

when "001010001001010" => rgb <= "100110";

when "001010001001011" => rgb <= "100110";

when "001010001001100" => rgb <= "100110";

when "001010001001101" => rgb <= "100110";

when "001010001001110" => rgb <= "100110";

when "001010001001111" => rgb <= "100110";

when "001010001010000" => rgb <= "000000";

when "001010101000111" => rgb <= "000000";

when "001010101001000" => rgb <= "100110";

when "001010101001001" => rgb <= "100110";

when "001010101001010" => rgb <= "100110";

when "001010101001011" => rgb <= "100110";

when "001010101001100" => rgb <= "100110";

when "001010101001101" => rgb <= "100110";

when "001010101001110" => rgb <= "100110";

when "001010101001111" => rgb <= "100110";

when "001010101010000" => rgb <= "000000";

when "001011001000111" => rgb <= "000000";

when "001011001001000" => rgb <= "100110";

when "001011001001001" => rgb <= "100110";

when "001011001001010" => rgb <= "100110";

when "001011001001011" => rgb <= "100110";

when "001011001001100" => rgb <= "100110";

when "001011001001101" => rgb <= "100110";

when "001011001001110" => rgb <= "100110";

when "001011001001111" => rgb <= "100110";

when "001011001010000" => rgb <= "000000";

when "001011101000111" => rgb <= "000000";

when "001011101001000" => rgb <= "100110";

when "001011101001001" => rgb <= "100110";

when "001011101001010" => rgb <= "100110";

when "001011101001011" => rgb <= "100110";

when "001011101001100" => rgb <= "100110";

when "001011101001101" => rgb <= "100110";

when "001011101001110" => rgb <= "100110";

when "001011101001111" => rgb <= "100110";

when "001011101010000" => rgb <= "000000";

when "001100001000111" => rgb <= "000000";

when "001100001001000" => rgb <= "100110";

when "001100001001001" => rgb <= "100110";

when "001100001001010" => rgb <= "100110";

when "001100001001011" => rgb <= "100110";

when "001100001001100" => rgb <= "100110";

when "001100001001101" => rgb <= "100110";

when "001100001001110" => rgb <= "100110";

when "001100001001111" => rgb <= "100110";

when "001100001010000" => rgb <= "000000";

when "001100101000111" => rgb <= "000000";

when "001100101001000" => rgb <= "100110";

when "001100101001001" => rgb <= "100110";

when "001100101001010" => rgb <= "100110";

when "001100101001011" => rgb <= "100110";

when "001100101001100" => rgb <= "100110";

when "001100101001101" => rgb <= "100110";

when "001100101001110" => rgb <= "100110";

when "001100101001111" => rgb <= "100110";

when "001100101010000" => rgb <= "000000";

when "001101001000111" => rgb <= "000000";

when "001101001001000" => rgb <= "100110";

when "001101001001001" => rgb <= "100110";

when "001101001001010" => rgb <= "100110";

when "001101001001011" => rgb <= "100110";

when "001101001001100" => rgb <= "100110";

when "001101001001101" => rgb <= "100110";

when "001101001001110" => rgb <= "100110";

when "001101001001111" => rgb <= "100110";

when "001101001010000" => rgb <= "000000";

when "001101101000111" => rgb <= "000000";

when "001101101001000" => rgb <= "100110";

when "001101101001001" => rgb <= "100110";

when "001101101001010" => rgb <= "100110";

when "001101101001011" => rgb <= "100110";

when "001101101001100" => rgb <= "100110";

when "001101101001101" => rgb <= "100110";

when "001101101001110" => rgb <= "100110";

when "001101101001111" => rgb <= "100110";

when "001101101010000" => rgb <= "000000";

when "001110001000111" => rgb <= "000000";

when "001110001001000" => rgb <= "100110";

when "001110001001001" => rgb <= "100110";

when "001110001001010" => rgb <= "100110";

when "001110001001011" => rgb <= "100110";

when "001110001001100" => rgb <= "100110";

when "001110001001101" => rgb <= "100110";

when "001110001001110" => rgb <= "100110";

when "001110001001111" => rgb <= "100110";

when "001110001010000" => rgb <= "000000";

when "001110101000111" => rgb <= "000000";

when "001110101001000" => rgb <= "100110";

when "001110101001001" => rgb <= "100110";

when "001110101001010" => rgb <= "100110";

when "001110101001011" => rgb <= "100110";

when "001110101001100" => rgb <= "100110";

when "001110101001101" => rgb <= "100110";

when "001110101001110" => rgb <= "100110";

when "001110101001111" => rgb <= "100110";

when "001110101010000" => rgb <= "000000";

when "001111001000111" => rgb <= "000000";

when "001111001001000" => rgb <= "100110";

when "001111001001001" => rgb <= "100110";

when "001111001001010" => rgb <= "100110";

when "001111001001011" => rgb <= "100110";

when "001111001001100" => rgb <= "100110";

when "001111001001101" => rgb <= "100110";

when "001111001001110" => rgb <= "100110";

when "001111001001111" => rgb <= "100110";

when "001111001010000" => rgb <= "000000";

when "001111101000111" => rgb <= "000000";

when "001111101001000" => rgb <= "100110";

when "001111101001001" => rgb <= "100110";

when "001111101001010" => rgb <= "100110";

when "001111101001011" => rgb <= "100110";

when "001111101001100" => rgb <= "100110";

when "001111101001101" => rgb <= "100110";

when "001111101001110" => rgb <= "100110";

when "001111101001111" => rgb <= "100110";

when "001111101010000" => rgb <= "000000";

when "010000001000111" => rgb <= "000000";

when "010000001001000" => rgb <= "100110";

when "010000001001001" => rgb <= "100110";

when "010000001001010" => rgb <= "100110";

when "010000001001011" => rgb <= "100110";

when "010000001001100" => rgb <= "100110";

when "010000001001101" => rgb <= "100110";

when "010000001001110" => rgb <= "100110";

when "010000001001111" => rgb <= "100110";

when "010000001010000" => rgb <= "000000";

when "010000101000111" => rgb <= "000000";

when "010000101001000" => rgb <= "100110";

when "010000101001001" => rgb <= "100110";

when "010000101001010" => rgb <= "100110";

when "010000101001011" => rgb <= "100110";

when "010000101001100" => rgb <= "100110";

when "010000101001101" => rgb <= "100110";

when "010000101001110" => rgb <= "100110";

when "010000101001111" => rgb <= "100110";

when "010000101010000" => rgb <= "000000";

when "010001001000111" => rgb <= "000000";

when "010001001001000" => rgb <= "100110";

when "010001001001001" => rgb <= "100110";

when "010001001001010" => rgb <= "100110";

when "010001001001011" => rgb <= "100110";

when "010001001001100" => rgb <= "100110";

when "010001001001101" => rgb <= "100110";

when "010001001001110" => rgb <= "100110";

when "010001001001111" => rgb <= "100110";

when "010001001010000" => rgb <= "000000";

when "010001101000111" => rgb <= "000000";

when "010001101001000" => rgb <= "100110";

when "010001101001001" => rgb <= "100110";

when "010001101001010" => rgb <= "100110";

when "010001101001011" => rgb <= "100110";

when "010001101001100" => rgb <= "100110";

when "010001101001101" => rgb <= "100110";

when "010001101001110" => rgb <= "100110";

when "010001101001111" => rgb <= "100110";

when "010001101010000" => rgb <= "000000";

when "010010001000111" => rgb <= "000000";

when "010010001001000" => rgb <= "100110";

when "010010001001001" => rgb <= "100110";

when "010010001001010" => rgb <= "100110";

when "010010001001011" => rgb <= "100110";

when "010010001001100" => rgb <= "100110";

when "010010001001101" => rgb <= "100110";

when "010010001001110" => rgb <= "100110";

when "010010001001111" => rgb <= "100110";

when "010010001010000" => rgb <= "000000";

when "010010101000111" => rgb <= "000000";

when "010010101001000" => rgb <= "100110";

when "010010101001001" => rgb <= "100110";

when "010010101001010" => rgb <= "100110";

when "010010101001011" => rgb <= "100110";

when "010010101001100" => rgb <= "100110";

when "010010101001101" => rgb <= "100110";

when "010010101001110" => rgb <= "100110";

when "010010101001111" => rgb <= "100110";

when "010010101010000" => rgb <= "000000";

when "010011001000111" => rgb <= "000000";

when "010011001001000" => rgb <= "100110";

when "010011001001001" => rgb <= "100110";

when "010011001001010" => rgb <= "100110";

when "010011001001011" => rgb <= "100110";

when "010011001001100" => rgb <= "100110";

when "010011001001101" => rgb <= "100110";

when "010011001001110" => rgb <= "100110";

when "010011001001111" => rgb <= "100110";

when "010011001010000" => rgb <= "000000";

when "010011101000111" => rgb <= "000000";

when "010011101001000" => rgb <= "100110";

when "010011101001001" => rgb <= "100110";

when "010011101001010" => rgb <= "100110";

when "010011101001011" => rgb <= "100110";

when "010011101001100" => rgb <= "100110";

when "010011101001101" => rgb <= "100110";

when "010011101001110" => rgb <= "100110";

when "010011101001111" => rgb <= "100110";

when "010011101010000" => rgb <= "000000";

when "010100001000111" => rgb <= "000000";

when "010100001001000" => rgb <= "100110";

when "010100001001001" => rgb <= "100110";

when "010100001001010" => rgb <= "100110";

when "010100001001011" => rgb <= "100110";

when "010100001001100" => rgb <= "100110";

when "010100001001101" => rgb <= "100110";

when "010100001001110" => rgb <= "100110";

when "010100001001111" => rgb <= "100110";

when "010100001010000" => rgb <= "000000";

when "010100101000111" => rgb <= "000000";

when "010100101001000" => rgb <= "100110";

when "010100101001001" => rgb <= "100110";

when "010100101001010" => rgb <= "100110";

when "010100101001011" => rgb <= "100110";

when "010100101001100" => rgb <= "100110";

when "010100101001101" => rgb <= "100110";

when "010100101001110" => rgb <= "100110";

when "010100101001111" => rgb <= "100110";

when "010100101010000" => rgb <= "000000";

when "010101001000111" => rgb <= "000000";

when "010101001001000" => rgb <= "100110";

when "010101001001001" => rgb <= "100110";

when "010101001001010" => rgb <= "100110";

when "010101001001011" => rgb <= "100110";

when "010101001001100" => rgb <= "100110";

when "010101001001101" => rgb <= "100110";

when "010101001001110" => rgb <= "100110";

when "010101001001111" => rgb <= "100110";

when "010101001010000" => rgb <= "000000";

when "010101101000111" => rgb <= "000000";

when "010101101001000" => rgb <= "100110";

when "010101101001001" => rgb <= "100110";

when "010101101001010" => rgb <= "100110";

when "010101101001011" => rgb <= "100110";

when "010101101001100" => rgb <= "100110";

when "010101101001101" => rgb <= "100110";

when "010101101001110" => rgb <= "100110";

when "010101101001111" => rgb <= "100110";

when "010101101010000" => rgb <= "000000";

when "010110001000111" => rgb <= "000000";

when "010110001001000" => rgb <= "100110";

when "010110001001001" => rgb <= "100110";

when "010110001001010" => rgb <= "100110";

when "010110001001011" => rgb <= "100110";

when "010110001001100" => rgb <= "100110";

when "010110001001101" => rgb <= "100110";

when "010110001001110" => rgb <= "100110";

when "010110001001111" => rgb <= "100110";

when "010110001010000" => rgb <= "000000";

when "010110101000111" => rgb <= "000000";

when "010110101001000" => rgb <= "100110";

when "010110101001001" => rgb <= "100110";

when "010110101001010" => rgb <= "100110";

when "010110101001011" => rgb <= "100110";

when "010110101001100" => rgb <= "100110";

when "010110101001101" => rgb <= "100110";

when "010110101001110" => rgb <= "100110";

when "010110101001111" => rgb <= "100110";

when "010110101010000" => rgb <= "000000";

when "010111001000111" => rgb <= "000000";

when "010111001001000" => rgb <= "100110";

when "010111001001001" => rgb <= "100110";

when "010111001001010" => rgb <= "100110";

when "010111001001011" => rgb <= "100110";

when "010111001001100" => rgb <= "100110";

when "010111001001101" => rgb <= "100110";

when "010111001001110" => rgb <= "100110";

when "010111001001111" => rgb <= "100110";

when "010111001010000" => rgb <= "000000";

when "010111101000111" => rgb <= "000000";

when "010111101001000" => rgb <= "100110";

when "010111101001001" => rgb <= "100110";

when "010111101001010" => rgb <= "100110";

when "010111101001011" => rgb <= "100110";

when "010111101001100" => rgb <= "100110";

when "010111101001101" => rgb <= "100110";

when "010111101001110" => rgb <= "100110";

when "010111101001111" => rgb <= "100110";

when "010111101010000" => rgb <= "000000";

when "011000001000111" => rgb <= "000000";

when "011000001001000" => rgb <= "100110";

when "011000001001001" => rgb <= "100110";

when "011000001001010" => rgb <= "100110";

when "011000001001011" => rgb <= "100110";

when "011000001001100" => rgb <= "100110";

when "011000001001101" => rgb <= "100110";

when "011000001001110" => rgb <= "100110";

when "011000001001111" => rgb <= "100110";

when "011000001010000" => rgb <= "000000";

when "011000101000111" => rgb <= "000000";

when "011000101001000" => rgb <= "100110";

when "011000101001001" => rgb <= "100110";

when "011000101001010" => rgb <= "100110";

when "011000101001011" => rgb <= "100110";

when "011000101001100" => rgb <= "100110";

when "011000101001101" => rgb <= "100110";

when "011000101001110" => rgb <= "100110";

when "011000101001111" => rgb <= "100110";

when "011000101010000" => rgb <= "000000";

when "011001001000111" => rgb <= "000000";

when "011001001001000" => rgb <= "100110";

when "011001001001001" => rgb <= "100110";

when "011001001001010" => rgb <= "100110";

when "011001001001011" => rgb <= "100110";

when "011001001001100" => rgb <= "100110";

when "011001001001101" => rgb <= "100110";

when "011001001001110" => rgb <= "100110";

when "011001001001111" => rgb <= "100110";

when "011001001010000" => rgb <= "000000";

when "011001101000111" => rgb <= "000000";

when "011001101001000" => rgb <= "100110";

when "011001101001001" => rgb <= "100110";

when "011001101001010" => rgb <= "100110";

when "011001101001011" => rgb <= "100110";

when "011001101001100" => rgb <= "100110";

when "011001101001101" => rgb <= "100110";

when "011001101001110" => rgb <= "100110";

when "011001101001111" => rgb <= "100110";

when "011001101010000" => rgb <= "000000";

when "011010001000111" => rgb <= "000000";

when "011010001001000" => rgb <= "100110";

when "011010001001001" => rgb <= "100110";

when "011010001001010" => rgb <= "100110";

when "011010001001011" => rgb <= "100110";

when "011010001001100" => rgb <= "100110";

when "011010001001101" => rgb <= "100110";

when "011010001001110" => rgb <= "100110";

when "011010001001111" => rgb <= "100110";

when "011010001010000" => rgb <= "000000";

when "011010101000111" => rgb <= "000000";

when "011010101001000" => rgb <= "100110";

when "011010101001001" => rgb <= "100110";

when "011010101001010" => rgb <= "100110";

when "011010101001011" => rgb <= "100110";

when "011010101001100" => rgb <= "100110";

when "011010101001101" => rgb <= "100110";

when "011010101001110" => rgb <= "100110";

when "011010101001111" => rgb <= "100110";

when "011010101010000" => rgb <= "000000";

when "011011001000111" => rgb <= "000000";

when "011011001001000" => rgb <= "100110";

when "011011001001001" => rgb <= "100110";

when "011011001001010" => rgb <= "100110";

when "011011001001011" => rgb <= "100110";

when "011011001001100" => rgb <= "100110";

when "011011001001101" => rgb <= "100110";

when "011011001001110" => rgb <= "100110";

when "011011001001111" => rgb <= "100110";

when "011011001010000" => rgb <= "000000";

when "011011101000111" => rgb <= "000000";

when "011011101001000" => rgb <= "100110";

when "011011101001001" => rgb <= "100110";

when "011011101001010" => rgb <= "100110";

when "011011101001011" => rgb <= "100110";

when "011011101001100" => rgb <= "100110";

when "011011101001101" => rgb <= "100110";

when "011011101001110" => rgb <= "100110";

when "011011101001111" => rgb <= "100110";

when "011011101010000" => rgb <= "000000";

when "011100001000111" => rgb <= "000000";

when "011100001001000" => rgb <= "100110";

when "011100001001001" => rgb <= "100110";

when "011100001001010" => rgb <= "100110";

when "011100001001011" => rgb <= "100110";

when "011100001001100" => rgb <= "100110";

when "011100001001101" => rgb <= "100110";

when "011100001001110" => rgb <= "100110";

when "011100001001111" => rgb <= "100110";

when "011100001010000" => rgb <= "000000";

when "011100101000111" => rgb <= "000000";

when "011100101001000" => rgb <= "100110";

when "011100101001001" => rgb <= "100110";

when "011100101001010" => rgb <= "100110";

when "011100101001011" => rgb <= "100110";

when "011100101001100" => rgb <= "100110";

when "011100101001101" => rgb <= "100110";

when "011100101001110" => rgb <= "100110";

when "011100101001111" => rgb <= "100110";

when "011100101010000" => rgb <= "000000";

when "011101001000111" => rgb <= "000000";

when "011101001001000" => rgb <= "100110";

when "011101001001001" => rgb <= "100110";

when "011101001001010" => rgb <= "100110";

when "011101001001011" => rgb <= "100110";

when "011101001001100" => rgb <= "100110";

when "011101001001101" => rgb <= "100110";

when "011101001001110" => rgb <= "100110";

when "011101001001111" => rgb <= "100110";

when "011101001010000" => rgb <= "000000";

when "011101101000111" => rgb <= "000000";

when "011101101001000" => rgb <= "100110";

when "011101101001001" => rgb <= "100110";

when "011101101001010" => rgb <= "100110";

when "011101101001011" => rgb <= "100110";

when "011101101001100" => rgb <= "100110";

when "011101101001101" => rgb <= "100110";

when "011101101001110" => rgb <= "100110";

when "011101101001111" => rgb <= "100110";

when "011101101010000" => rgb <= "000000";

when "011110001000111" => rgb <= "000000";

when "011110001001000" => rgb <= "100110";

when "011110001001001" => rgb <= "100110";

when "011110001001010" => rgb <= "100110";

when "011110001001011" => rgb <= "100110";

when "011110001001100" => rgb <= "100110";

when "011110001001101" => rgb <= "100110";

when "011110001001110" => rgb <= "100110";

when "011110001001111" => rgb <= "100110";

when "011110001010000" => rgb <= "000000";

when "011110101000111" => rgb <= "000000";

when "011110101001000" => rgb <= "100110";

when "011110101001001" => rgb <= "100110";

when "011110101001010" => rgb <= "100110";

when "011110101001011" => rgb <= "100110";

when "011110101001100" => rgb <= "100110";

when "011110101001101" => rgb <= "100110";

when "011110101001110" => rgb <= "100110";

when "011110101001111" => rgb <= "100110";

when "011110101010000" => rgb <= "000000";

when "011111001000111" => rgb <= "000000";

when "011111001001000" => rgb <= "100110";

when "011111001001001" => rgb <= "100110";

when "011111001001010" => rgb <= "100110";

when "011111001001011" => rgb <= "100110";

when "011111001001100" => rgb <= "100110";

when "011111001001101" => rgb <= "100110";

when "011111001001110" => rgb <= "100110";

when "011111001001111" => rgb <= "100110";

when "011111001010000" => rgb <= "000000";

when "011111101000111" => rgb <= "000000";

when "011111101001000" => rgb <= "000000";

when "011111101001001" => rgb <= "000000";

when "011111101001010" => rgb <= "000000";

when "011111101001011" => rgb <= "000000";

when "011111101001100" => rgb <= "000000";

when "011111101001101" => rgb <= "000000";

when "011111101001110" => rgb <= "000000";

when "011111101001111" => rgb <= "000000";

when "011111101010000" => rgb <= "000000";
when others => rgb <= "111111"; --will update l8r
end case;
end if;
end process;
	addressOut <= address;
end;