library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;


entity startScreen is --rom for the background
port(
    clk : in std_logic;
	address : in unsigned (14 downto 0); 
    rgb : out unsigned(5 downto 0)
);
end startScreen;


architecture synth of startScreen is 

signal addressOut : unsigned(14 downto 0); 

begin
    process (clk) is begin
        if rising_edge(clk) then
            case addressOut is
			when "000101000010000" => rgb <= "000000";
when "000101000010001" => rgb <= "000000";
when "000101000010010" => rgb <= "000000";
when "000101000010011" => rgb <= "000000";
when "000101000010100" => rgb <= "000000";
when "000101000010101" => rgb <= "000000";
when "000101000010110" => rgb <= "000000";
when "000101000010111" => rgb <= "000000";
when "000101000011000" => rgb <= "000000";
when "000101000011001" => rgb <= "000000";
when "000101000011100" => rgb <= "000000";
when "000101000011101" => rgb <= "000000";
when "000101000011110" => rgb <= "000000";
when "000101000011111" => rgb <= "000000";
when "000101000100000" => rgb <= "000000";
when "000101000100001" => rgb <= "000000";
when "000101000100010" => rgb <= "000000";
when "000101000100011" => rgb <= "000000";
when "000101000100100" => rgb <= "000000";
when "000101000100101" => rgb <= "000000";
when "000101000100110" => rgb <= "000000";
when "000101000100111" => rgb <= "000000";
when "000101000101000" => rgb <= "000000";
when "000101000101001" => rgb <= "000000";
when "000101000101100" => rgb <= "000000";
when "000101000101101" => rgb <= "000000";
when "000101000101110" => rgb <= "000000";
when "000101000101111" => rgb <= "000000";
when "000101000110000" => rgb <= "000000";
when "000101000110001" => rgb <= "000000";
when "000101000110010" => rgb <= "000000";
when "000101000110011" => rgb <= "000000";
when "000101000110111" => rgb <= "000000";
when "000101000111000" => rgb <= "000000";
when "000101000111001" => rgb <= "000000";
when "000101000111010" => rgb <= "000000";
when "000101000111011" => rgb <= "000000";
when "000101000111100" => rgb <= "000000";
when "000101000111101" => rgb <= "000000";
when "000101000111110" => rgb <= "000000";
when "000101000111111" => rgb <= "000000";
when "000101001000000" => rgb <= "000000";
when "000101001000001" => rgb <= "000000";
when "000101001000010" => rgb <= "000000";
when "000101001000100" => rgb <= "000000";
when "000101001000101" => rgb <= "000000";
when "000101001000110" => rgb <= "000000";
when "000101001000111" => rgb <= "000000";
when "000101001001000" => rgb <= "000000";
when "000101001001001" => rgb <= "000000";
when "000101001001010" => rgb <= "000000";
when "000101001001011" => rgb <= "000000";
when "000101001001100" => rgb <= "000000";
when "000101001001101" => rgb <= "000000";
when "000101001001110" => rgb <= "000000";
when "000101001001111" => rgb <= "000000";
when "000101001010000" => rgb <= "000000";
when "000101001011100" => rgb <= "000000";
when "000101001011101" => rgb <= "000000";
when "000101001011110" => rgb <= "000000";
when "000101001011111" => rgb <= "000000";
when "000101001100000" => rgb <= "000000";
when "000101001100001" => rgb <= "000000";
when "000101001100010" => rgb <= "000000";
when "000101001100011" => rgb <= "000000";
when "000101001100100" => rgb <= "000000";
when "000101001100101" => rgb <= "000000";
when "000101001101010" => rgb <= "000000";
when "000101001101011" => rgb <= "000000";
when "000101001101100" => rgb <= "000000";
when "000101001101101" => rgb <= "000000";
when "000101001101110" => rgb <= "000000";
when "000101001101111" => rgb <= "000000";
when "000101001110000" => rgb <= "000000";
when "000101001110001" => rgb <= "000000";
when "000101001110101" => rgb <= "000000";
when "000101001110110" => rgb <= "000000";
when "000101001110111" => rgb <= "000000";
when "000101001111000" => rgb <= "000000";
when "000101001111001" => rgb <= "000000";
when "000101001111010" => rgb <= "000000";
when "000101001111110" => rgb <= "000000";
when "000101001111111" => rgb <= "000000";
when "000101010000000" => rgb <= "000000";
when "000101010000001" => rgb <= "000000";
when "000101010000010" => rgb <= "000000";
when "000101010000011" => rgb <= "000000";
when "000101010000100" => rgb <= "000000";
when "000101010000101" => rgb <= "000000";
when "000101010000110" => rgb <= "000000";
when "000101010000111" => rgb <= "000000";
when "000101010001000" => rgb <= "000000";
when "000101010001001" => rgb <= "000000";
when "000101010001010" => rgb <= "000000";
when "000101010001011" => rgb <= "000000";
when "000101010001100" => rgb <= "000000";
when "000101010001101" => rgb <= "000000";
when "000101010001110" => rgb <= "000000";
when "000101010001111" => rgb <= "000000";
when "000101100010000" => rgb <= "000000";
when "000101100010001" => rgb <= "100110";
when "000101100010010" => rgb <= "100110";
when "000101100010011" => rgb <= "100110";
when "000101100010100" => rgb <= "100110";
when "000101100010101" => rgb <= "100110";
when "000101100010110" => rgb <= "100110";
when "000101100010111" => rgb <= "100110";
when "000101100011000" => rgb <= "100110";
when "000101100011001" => rgb <= "000000";
when "000101100011010" => rgb <= "000000";
when "000101100011011" => rgb <= "000000";
when "000101100011100" => rgb <= "000000";
when "000101100011101" => rgb <= "100110";
when "000101100011110" => rgb <= "100110";
when "000101100011111" => rgb <= "100110";
when "000101100100000" => rgb <= "100110";
when "000101100100001" => rgb <= "100110";
when "000101100100010" => rgb <= "100110";
when "000101100100011" => rgb <= "100110";
when "000101100100100" => rgb <= "100110";
when "000101100100101" => rgb <= "100110";
when "000101100100110" => rgb <= "100110";
when "000101100100111" => rgb <= "100110";
when "000101100101000" => rgb <= "000000";
when "000101100101001" => rgb <= "000000";
when "000101100101010" => rgb <= "000000";
when "000101100101011" => rgb <= "000000";
when "000101100101100" => rgb <= "000000";
when "000101100101101" => rgb <= "100110";
when "000101100101110" => rgb <= "100110";
when "000101100101111" => rgb <= "100110";
when "000101100110000" => rgb <= "100110";
when "000101100110001" => rgb <= "100110";
when "000101100110010" => rgb <= "100110";
when "000101100110011" => rgb <= "000000";
when "000101100110100" => rgb <= "000000";
when "000101100110101" => rgb <= "000000";
when "000101100110111" => rgb <= "000000";
when "000101100111000" => rgb <= "100110";
when "000101100111001" => rgb <= "100110";
when "000101100111010" => rgb <= "100110";
when "000101100111011" => rgb <= "100110";
when "000101100111100" => rgb <= "100110";
when "000101100111101" => rgb <= "100110";
when "000101100111110" => rgb <= "100110";
when "000101100111111" => rgb <= "100110";
when "000101101000000" => rgb <= "100110";
when "000101101000001" => rgb <= "000000";
when "000101101000010" => rgb <= "000000";
when "000101101000011" => rgb <= "000000";
when "000101101000100" => rgb <= "000000";
when "000101101000101" => rgb <= "100110";
when "000101101000110" => rgb <= "100110";
when "000101101000111" => rgb <= "100110";
when "000101101001000" => rgb <= "100110";
when "000101101001001" => rgb <= "100110";
when "000101101001010" => rgb <= "100110";
when "000101101001011" => rgb <= "100110";
when "000101101001100" => rgb <= "100110";
when "000101101001101" => rgb <= "100110";
when "000101101001110" => rgb <= "100110";
when "000101101001111" => rgb <= "100110";
when "000101101010000" => rgb <= "000000";
when "000101101010001" => rgb <= "000000";
when "000101101010010" => rgb <= "000000";
when "000101101011010" => rgb <= "000000";
when "000101101011011" => rgb <= "000000";
when "000101101011100" => rgb <= "000000";
when "000101101011101" => rgb <= "100110";
when "000101101011110" => rgb <= "100110";
when "000101101011111" => rgb <= "100110";
when "000101101100000" => rgb <= "100110";
when "000101101100001" => rgb <= "100110";
when "000101101100010" => rgb <= "100110";
when "000101101100011" => rgb <= "100110";
when "000101101100100" => rgb <= "100110";
when "000101101100101" => rgb <= "000000";
when "000101101100110" => rgb <= "000000";
when "000101101101010" => rgb <= "000000";
when "000101101101011" => rgb <= "100110";
when "000101101101100" => rgb <= "100110";
when "000101101101101" => rgb <= "100110";
when "000101101101110" => rgb <= "100110";
when "000101101101111" => rgb <= "100110";
when "000101101110000" => rgb <= "100110";
when "000101101110001" => rgb <= "000000";
when "000101101110010" => rgb <= "000000";
when "000101101110011" => rgb <= "000000";
when "000101101110101" => rgb <= "000000";
when "000101101110110" => rgb <= "100110";
when "000101101110111" => rgb <= "100110";
when "000101101111000" => rgb <= "100110";
when "000101101111001" => rgb <= "100110";
when "000101101111010" => rgb <= "000000";
when "000101101111011" => rgb <= "000000";
when "000101101111110" => rgb <= "000000";
when "000101101111111" => rgb <= "100110";
when "000101110000000" => rgb <= "100110";
when "000101110000001" => rgb <= "100110";
when "000101110000010" => rgb <= "100110";
when "000101110000011" => rgb <= "000000";
when "000101110000100" => rgb <= "000000";
when "000101110000101" => rgb <= "100110";
when "000101110000110" => rgb <= "100110";
when "000101110000111" => rgb <= "100110";
when "000101110001000" => rgb <= "100110";
when "000101110001001" => rgb <= "100110";
when "000101110001010" => rgb <= "100110";
when "000101110001011" => rgb <= "100110";
when "000101110001100" => rgb <= "100110";
when "000101110001101" => rgb <= "100110";
when "000101110001110" => rgb <= "100110";
when "000101110001111" => rgb <= "000000";
when "000101110010000" => rgb <= "000000";
when "000101110010001" => rgb <= "000000";
when "000110000001110" => rgb <= "000000";
when "000110000001111" => rgb <= "000000";
when "000110000010000" => rgb <= "000000";
when "000110000010001" => rgb <= "100110";
when "000110000010010" => rgb <= "100110";
when "000110000010011" => rgb <= "100110";
when "000110000010100" => rgb <= "100110";
when "000110000010101" => rgb <= "100110";
when "000110000010110" => rgb <= "100110";
when "000110000010111" => rgb <= "100110";
when "000110000011000" => rgb <= "100110";
when "000110000011001" => rgb <= "000000";
when "000110000011010" => rgb <= "000000";
when "000110000011011" => rgb <= "000000";
when "000110000011100" => rgb <= "000000";
when "000110000011101" => rgb <= "100110";
when "000110000011110" => rgb <= "100110";
when "000110000011111" => rgb <= "100110";
when "000110000100000" => rgb <= "100110";
when "000110000100001" => rgb <= "100110";
when "000110000100010" => rgb <= "100110";
when "000110000100011" => rgb <= "100110";
when "000110000100100" => rgb <= "100110";
when "000110000100101" => rgb <= "100110";
when "000110000100110" => rgb <= "100110";
when "000110000100111" => rgb <= "100110";
when "000110000101000" => rgb <= "000000";
when "000110000101001" => rgb <= "000000";
when "000110000101010" => rgb <= "000000";
when "000110000101011" => rgb <= "000000";
when "000110000101100" => rgb <= "000000";
when "000110000101101" => rgb <= "100110";
when "000110000101110" => rgb <= "100110";
when "000110000101111" => rgb <= "100110";
when "000110000110000" => rgb <= "100110";
when "000110000110001" => rgb <= "100110";
when "000110000110010" => rgb <= "100110";
when "000110000110011" => rgb <= "000000";
when "000110000110100" => rgb <= "000000";
when "000110000110101" => rgb <= "000000";
when "000110000110110" => rgb <= "000000";
when "000110000110111" => rgb <= "000000";
when "000110000111000" => rgb <= "100110";
when "000110000111001" => rgb <= "100110";
when "000110000111010" => rgb <= "100110";
when "000110000111011" => rgb <= "100110";
when "000110000111100" => rgb <= "100110";
when "000110000111101" => rgb <= "100110";
when "000110000111110" => rgb <= "100110";
when "000110000111111" => rgb <= "100110";
when "000110001000000" => rgb <= "100110";
when "000110001000001" => rgb <= "100110";
when "000110001000010" => rgb <= "100110";
when "000110001000011" => rgb <= "000000";
when "000110001000100" => rgb <= "000000";
when "000110001000101" => rgb <= "100110";
when "000110001000110" => rgb <= "100110";
when "000110001000111" => rgb <= "100110";
when "000110001001000" => rgb <= "100110";
when "000110001001001" => rgb <= "100110";
when "000110001001010" => rgb <= "100110";
when "000110001001011" => rgb <= "100110";
when "000110001001100" => rgb <= "100110";
when "000110001001101" => rgb <= "100110";
when "000110001001110" => rgb <= "100110";
when "000110001001111" => rgb <= "100110";
when "000110001010000" => rgb <= "000000";
when "000110001010001" => rgb <= "000000";
when "000110001010010" => rgb <= "000000";
when "000110001011001" => rgb <= "000000";
when "000110001011010" => rgb <= "000000";
when "000110001011011" => rgb <= "100110";
when "000110001011100" => rgb <= "100110";
when "000110001011101" => rgb <= "100110";
when "000110001011110" => rgb <= "100110";
when "000110001011111" => rgb <= "100110";
when "000110001100000" => rgb <= "100110";
when "000110001100001" => rgb <= "100110";
when "000110001100010" => rgb <= "100110";
when "000110001100011" => rgb <= "100110";
when "000110001100100" => rgb <= "100110";
when "000110001100101" => rgb <= "100110";
when "000110001100110" => rgb <= "000000";
when "000110001100111" => rgb <= "000000";
when "000110001101000" => rgb <= "000000";
when "000110001101001" => rgb <= "000000";
when "000110001101010" => rgb <= "000000";
when "000110001101011" => rgb <= "100110";
when "000110001101100" => rgb <= "100110";
when "000110001101101" => rgb <= "100110";
when "000110001101110" => rgb <= "100110";
when "000110001101111" => rgb <= "100110";
when "000110001110000" => rgb <= "100110";
when "000110001110001" => rgb <= "000000";
when "000110001110010" => rgb <= "000000";
when "000110001110011" => rgb <= "000000";
when "000110001110100" => rgb <= "000000";
when "000110001110101" => rgb <= "000000";
when "000110001110110" => rgb <= "100110";
when "000110001110111" => rgb <= "100110";
when "000110001111000" => rgb <= "100110";
when "000110001111001" => rgb <= "100110";
when "000110001111010" => rgb <= "000000";
when "000110001111011" => rgb <= "000000";
when "000110001111100" => rgb <= "000000";
when "000110001111101" => rgb <= "000000";
when "000110001111110" => rgb <= "000000";
when "000110001111111" => rgb <= "100110";
when "000110010000000" => rgb <= "100110";
when "000110010000001" => rgb <= "100110";
when "000110010000010" => rgb <= "100110";
when "000110010000011" => rgb <= "000000";
when "000110010000100" => rgb <= "000000";
when "000110010000101" => rgb <= "100110";
when "000110010000110" => rgb <= "100110";
when "000110010000111" => rgb <= "100110";
when "000110010001000" => rgb <= "100110";
when "000110010001001" => rgb <= "100110";
when "000110010001010" => rgb <= "100110";
when "000110010001011" => rgb <= "100110";
when "000110010001100" => rgb <= "100110";
when "000110010001101" => rgb <= "100110";
when "000110010001110" => rgb <= "100110";
when "000110010001111" => rgb <= "000000";
when "000110010010000" => rgb <= "000000";
when "000110010010001" => rgb <= "000000";
when "000110100001110" => rgb <= "000000";
when "000110100001111" => rgb <= "100110";
when "000110100010000" => rgb <= "100110";
when "000110100010001" => rgb <= "100110";
when "000110100010010" => rgb <= "100110";
when "000110100010011" => rgb <= "100110";
when "000110100010100" => rgb <= "100110";
when "000110100010101" => rgb <= "100110";
when "000110100010110" => rgb <= "100110";
when "000110100010111" => rgb <= "100110";
when "000110100011000" => rgb <= "100110";
when "000110100011001" => rgb <= "100110";
when "000110100011010" => rgb <= "100110";
when "000110100011011" => rgb <= "000000";
when "000110100011100" => rgb <= "000000";
when "000110100011101" => rgb <= "100110";
when "000110100011110" => rgb <= "100110";
when "000110100011111" => rgb <= "100110";
when "000110100100000" => rgb <= "100110";
when "000110100100001" => rgb <= "100110";
when "000110100100010" => rgb <= "100110";
when "000110100100011" => rgb <= "100110";
when "000110100100100" => rgb <= "100110";
when "000110100100101" => rgb <= "100110";
when "000110100100110" => rgb <= "100110";
when "000110100100111" => rgb <= "100110";
when "000110100101000" => rgb <= "000000";
when "000110100101001" => rgb <= "000000";
when "000110100101010" => rgb <= "000000";
when "000110100101011" => rgb <= "100110";
when "000110100101100" => rgb <= "100110";
when "000110100101101" => rgb <= "100110";
when "000110100101110" => rgb <= "100110";
when "000110100101111" => rgb <= "100110";
when "000110100110000" => rgb <= "100110";
when "000110100110001" => rgb <= "100110";
when "000110100110010" => rgb <= "100110";
when "000110100110011" => rgb <= "100110";
when "000110100110100" => rgb <= "100110";
when "000110100110101" => rgb <= "000000";
when "000110100110110" => rgb <= "000000";
when "000110100110111" => rgb <= "000000";
when "000110100111000" => rgb <= "100110";
when "000110100111001" => rgb <= "100110";
when "000110100111010" => rgb <= "100110";
when "000110100111011" => rgb <= "000000";
when "000110100111100" => rgb <= "000000";
when "000110100111101" => rgb <= "000000";
when "000110100111110" => rgb <= "000000";
when "000110100111111" => rgb <= "000000";
when "000110101000000" => rgb <= "100110";
when "000110101000001" => rgb <= "100110";
when "000110101000010" => rgb <= "100110";
when "000110101000011" => rgb <= "000000";
when "000110101000100" => rgb <= "000000";
when "000110101000101" => rgb <= "100110";
when "000110101000110" => rgb <= "100110";
when "000110101000111" => rgb <= "100110";
when "000110101001000" => rgb <= "100110";
when "000110101001001" => rgb <= "100110";
when "000110101001010" => rgb <= "100110";
when "000110101001011" => rgb <= "100110";
when "000110101001100" => rgb <= "100110";
when "000110101001101" => rgb <= "100110";
when "000110101001110" => rgb <= "100110";
when "000110101001111" => rgb <= "100110";
when "000110101010000" => rgb <= "000000";
when "000110101010001" => rgb <= "000000";
when "000110101010010" => rgb <= "000000";
when "000110101011001" => rgb <= "000000";
when "000110101011010" => rgb <= "100110";
when "000110101011011" => rgb <= "100110";
when "000110101011100" => rgb <= "100110";
when "000110101011101" => rgb <= "100110";
when "000110101011110" => rgb <= "100110";
when "000110101011111" => rgb <= "100110";
when "000110101100000" => rgb <= "100110";
when "000110101100001" => rgb <= "100110";
when "000110101100010" => rgb <= "100110";
when "000110101100011" => rgb <= "100110";
when "000110101100100" => rgb <= "100110";
when "000110101100101" => rgb <= "100110";
when "000110101100110" => rgb <= "000000";
when "000110101100111" => rgb <= "000000";
when "000110101101000" => rgb <= "000000";
when "000110101101001" => rgb <= "100110";
when "000110101101010" => rgb <= "100110";
when "000110101101011" => rgb <= "100110";
when "000110101101100" => rgb <= "100110";
when "000110101101101" => rgb <= "100110";
when "000110101101110" => rgb <= "100110";
when "000110101101111" => rgb <= "100110";
when "000110101110000" => rgb <= "100110";
when "000110101110001" => rgb <= "100110";
when "000110101110010" => rgb <= "100110";
when "000110101110011" => rgb <= "000000";
when "000110101110100" => rgb <= "000000";
when "000110101110101" => rgb <= "000000";
when "000110101110110" => rgb <= "100110";
when "000110101110111" => rgb <= "100110";
when "000110101111000" => rgb <= "100110";
when "000110101111001" => rgb <= "100110";
when "000110101111010" => rgb <= "100110";
when "000110101111011" => rgb <= "000000";
when "000110101111100" => rgb <= "000000";
when "000110101111101" => rgb <= "000000";
when "000110101111110" => rgb <= "100110";
when "000110101111111" => rgb <= "100110";
when "000110110000000" => rgb <= "100110";
when "000110110000001" => rgb <= "100110";
when "000110110000010" => rgb <= "100110";
when "000110110000011" => rgb <= "000000";
when "000110110000100" => rgb <= "000000";
when "000110110000101" => rgb <= "100110";
when "000110110000110" => rgb <= "100110";
when "000110110000111" => rgb <= "100110";
when "000110110001000" => rgb <= "100110";
when "000110110001001" => rgb <= "100110";
when "000110110001010" => rgb <= "100110";
when "000110110001011" => rgb <= "100110";
when "000110110001100" => rgb <= "100110";
when "000110110001101" => rgb <= "100110";
when "000110110001110" => rgb <= "100110";
when "000110110001111" => rgb <= "000000";
when "000110110010000" => rgb <= "000000";
when "000110110010001" => rgb <= "000000";
when "000111000001110" => rgb <= "000000";
when "000111000001111" => rgb <= "100110";
when "000111000010000" => rgb <= "100110";
when "000111000010001" => rgb <= "100110";
when "000111000010010" => rgb <= "100110";
when "000111000010011" => rgb <= "000000";
when "000111000010100" => rgb <= "000000";
when "000111000010101" => rgb <= "000000";
when "000111000010110" => rgb <= "000000";
when "000111000010111" => rgb <= "100110";
when "000111000011000" => rgb <= "100110";
when "000111000011001" => rgb <= "100110";
when "000111000011010" => rgb <= "100110";
when "000111000011011" => rgb <= "000000";
when "000111000011100" => rgb <= "000000";
when "000111000011101" => rgb <= "000000";
when "000111000011110" => rgb <= "000000";
when "000111000011111" => rgb <= "000000";
when "000111000100000" => rgb <= "000000";
when "000111000100001" => rgb <= "100110";
when "000111000100010" => rgb <= "100110";
when "000111000100011" => rgb <= "100110";
when "000111000100100" => rgb <= "000000";
when "000111000100101" => rgb <= "000000";
when "000111000100110" => rgb <= "000000";
when "000111000100111" => rgb <= "000000";
when "000111000101000" => rgb <= "000000";
when "000111000101001" => rgb <= "000000";
when "000111000101010" => rgb <= "000000";
when "000111000101011" => rgb <= "100110";
when "000111000101100" => rgb <= "100110";
when "000111000101101" => rgb <= "100110";
when "000111000101110" => rgb <= "000000";
when "000111000101111" => rgb <= "000000";
when "000111000110000" => rgb <= "000000";
when "000111000110001" => rgb <= "000000";
when "000111000110010" => rgb <= "100110";
when "000111000110011" => rgb <= "100110";
when "000111000110100" => rgb <= "100110";
when "000111000110101" => rgb <= "000000";
when "000111000110110" => rgb <= "000000";
when "000111000110111" => rgb <= "000000";
when "000111000111000" => rgb <= "100110";
when "000111000111001" => rgb <= "100110";
when "000111000111010" => rgb <= "100110";
when "000111000111011" => rgb <= "000000";
when "000111000111100" => rgb <= "000000";
when "000111000111101" => rgb <= "000000";
when "000111000111110" => rgb <= "000000";
when "000111000111111" => rgb <= "000000";
when "000111001000000" => rgb <= "100110";
when "000111001000001" => rgb <= "100110";
when "000111001000010" => rgb <= "100110";
when "000111001000011" => rgb <= "000000";
when "000111001000100" => rgb <= "000000";
when "000111001000101" => rgb <= "000000";
when "000111001000110" => rgb <= "000000";
when "000111001000111" => rgb <= "000000";
when "000111001001000" => rgb <= "000000";
when "000111001001001" => rgb <= "100110";
when "000111001001010" => rgb <= "100110";
when "000111001001011" => rgb <= "100110";
when "000111001001100" => rgb <= "000000";
when "000111001001101" => rgb <= "000000";
when "000111001001110" => rgb <= "000000";
when "000111001001111" => rgb <= "000000";
when "000111001010000" => rgb <= "000000";
when "000111001010001" => rgb <= "000000";
when "000111001010010" => rgb <= "000000";
when "000111001011001" => rgb <= "000000";
when "000111001011010" => rgb <= "100110";
when "000111001011011" => rgb <= "100110";
when "000111001011100" => rgb <= "100110";
when "000111001011101" => rgb <= "100110";
when "000111001011110" => rgb <= "000000";
when "000111001011111" => rgb <= "000000";
when "000111001100000" => rgb <= "000000";
when "000111001100001" => rgb <= "000000";
when "000111001100010" => rgb <= "000000";
when "000111001100011" => rgb <= "100110";
when "000111001100100" => rgb <= "100110";
when "000111001100101" => rgb <= "100110";
when "000111001100110" => rgb <= "000000";
when "000111001100111" => rgb <= "000000";
when "000111001101000" => rgb <= "000000";
when "000111001101001" => rgb <= "100110";
when "000111001101010" => rgb <= "100110";
when "000111001101011" => rgb <= "100110";
when "000111001101100" => rgb <= "000000";
when "000111001101101" => rgb <= "000000";
when "000111001101110" => rgb <= "000000";
when "000111001101111" => rgb <= "000000";
when "000111001110000" => rgb <= "100110";
when "000111001110001" => rgb <= "100110";
when "000111001110010" => rgb <= "100110";
when "000111001110011" => rgb <= "000000";
when "000111001110100" => rgb <= "000000";
when "000111001110101" => rgb <= "000000";
when "000111001110110" => rgb <= "100110";
when "000111001110111" => rgb <= "100110";
when "000111001111000" => rgb <= "100110";
when "000111001111001" => rgb <= "100110";
when "000111001111010" => rgb <= "100110";
when "000111001111011" => rgb <= "000000";
when "000111001111100" => rgb <= "000000";
when "000111001111101" => rgb <= "000000";
when "000111001111110" => rgb <= "100110";
when "000111001111111" => rgb <= "100110";
when "000111010000000" => rgb <= "100110";
when "000111010000001" => rgb <= "100110";
when "000111010000010" => rgb <= "100110";
when "000111010000011" => rgb <= "000000";
when "000111010000100" => rgb <= "000000";
when "000111010000101" => rgb <= "100110";
when "000111010000110" => rgb <= "100110";
when "000111010000111" => rgb <= "100110";
when "000111010001000" => rgb <= "000000";
when "000111010001001" => rgb <= "000000";
when "000111010001010" => rgb <= "000000";
when "000111010001011" => rgb <= "000000";
when "000111010001100" => rgb <= "000000";
when "000111010001101" => rgb <= "000000";
when "000111010001110" => rgb <= "000000";
when "000111010001111" => rgb <= "000000";
when "000111010010000" => rgb <= "000000";
when "000111010010001" => rgb <= "000000";
when "000111100001110" => rgb <= "000000";
when "000111100001111" => rgb <= "100110";
when "000111100010000" => rgb <= "100110";
when "000111100010001" => rgb <= "100110";
when "000111100010010" => rgb <= "100110";
when "000111100010011" => rgb <= "000000";
when "000111100010100" => rgb <= "000000";
when "000111100010101" => rgb <= "000000";
when "000111100010110" => rgb <= "000000";
when "000111100010111" => rgb <= "100110";
when "000111100011000" => rgb <= "100110";
when "000111100011001" => rgb <= "100110";
when "000111100011010" => rgb <= "100110";
when "000111100011011" => rgb <= "000000";
when "000111100011100" => rgb <= "000000";
when "000111100011101" => rgb <= "000000";
when "000111100011110" => rgb <= "000000";
when "000111100011111" => rgb <= "000000";
when "000111100100000" => rgb <= "000000";
when "000111100100001" => rgb <= "100110";
when "000111100100010" => rgb <= "100110";
when "000111100100011" => rgb <= "100110";
when "000111100100100" => rgb <= "000000";
when "000111100100101" => rgb <= "000000";
when "000111100100110" => rgb <= "000000";
when "000111100100111" => rgb <= "000000";
when "000111100101000" => rgb <= "000000";
when "000111100101001" => rgb <= "000000";
when "000111100101010" => rgb <= "000000";
when "000111100101011" => rgb <= "100110";
when "000111100101100" => rgb <= "100110";
when "000111100101101" => rgb <= "100110";
when "000111100101110" => rgb <= "000000";
when "000111100101111" => rgb <= "000000";
when "000111100110000" => rgb <= "000000";
when "000111100110001" => rgb <= "000000";
when "000111100110010" => rgb <= "100110";
when "000111100110011" => rgb <= "100110";
when "000111100110100" => rgb <= "100110";
when "000111100110101" => rgb <= "000000";
when "000111100110110" => rgb <= "000000";
when "000111100110111" => rgb <= "000000";
when "000111100111000" => rgb <= "100110";
when "000111100111001" => rgb <= "100110";
when "000111100111010" => rgb <= "100110";
when "000111100111011" => rgb <= "000000";
when "000111100111100" => rgb <= "000000";
when "000111100111101" => rgb <= "000000";
when "000111100111110" => rgb <= "000000";
when "000111100111111" => rgb <= "000000";
when "000111101000000" => rgb <= "100110";
when "000111101000001" => rgb <= "100110";
when "000111101000010" => rgb <= "100110";
when "000111101000011" => rgb <= "000000";
when "000111101000100" => rgb <= "000000";
when "000111101000101" => rgb <= "000000";
when "000111101000110" => rgb <= "000000";
when "000111101000111" => rgb <= "000000";
when "000111101001000" => rgb <= "000000";
when "000111101001001" => rgb <= "100110";
when "000111101001010" => rgb <= "100110";
when "000111101001011" => rgb <= "100110";
when "000111101001100" => rgb <= "000000";
when "000111101001101" => rgb <= "000000";
when "000111101001110" => rgb <= "000000";
when "000111101001111" => rgb <= "000000";
when "000111101010000" => rgb <= "000000";
when "000111101010001" => rgb <= "000000";
when "000111101010010" => rgb <= "000000";
when "000111101011001" => rgb <= "000000";
when "000111101011010" => rgb <= "100110";
when "000111101011011" => rgb <= "100110";
when "000111101011100" => rgb <= "100110";
when "000111101011101" => rgb <= "000000";
when "000111101011110" => rgb <= "000000";
when "000111101011111" => rgb <= "000000";
when "000111101100000" => rgb <= "000000";
when "000111101100001" => rgb <= "000000";
when "000111101100010" => rgb <= "000000";
when "000111101100011" => rgb <= "000000";
when "000111101100100" => rgb <= "000000";
when "000111101100101" => rgb <= "000000";
when "000111101100110" => rgb <= "000000";
when "000111101100111" => rgb <= "000000";
when "000111101101000" => rgb <= "000000";
when "000111101101001" => rgb <= "100110";
when "000111101101010" => rgb <= "100110";
when "000111101101011" => rgb <= "100110";
when "000111101101100" => rgb <= "000000";
when "000111101101101" => rgb <= "000000";
when "000111101101110" => rgb <= "000000";
when "000111101101111" => rgb <= "000000";
when "000111101110000" => rgb <= "100110";
when "000111101110001" => rgb <= "100110";
when "000111101110010" => rgb <= "100110";
when "000111101110011" => rgb <= "000000";
when "000111101110100" => rgb <= "000000";
when "000111101110101" => rgb <= "000000";
when "000111101110110" => rgb <= "100110";
when "000111101110111" => rgb <= "100110";
when "000111101111000" => rgb <= "100110";
when "000111101111001" => rgb <= "100110";
when "000111101111010" => rgb <= "100110";
when "000111101111011" => rgb <= "100110";
when "000111101111100" => rgb <= "000000";
when "000111101111101" => rgb <= "100110";
when "000111101111110" => rgb <= "100110";
when "000111101111111" => rgb <= "100110";
when "000111110000000" => rgb <= "100110";
when "000111110000001" => rgb <= "100110";
when "000111110000010" => rgb <= "100110";
when "000111110000011" => rgb <= "000000";
when "000111110000100" => rgb <= "000000";
when "000111110000101" => rgb <= "100110";
when "000111110000110" => rgb <= "100110";
when "000111110000111" => rgb <= "100110";
when "000111110001000" => rgb <= "000000";
when "000111110001001" => rgb <= "000000";
when "000111110001010" => rgb <= "000000";
when "000111110001011" => rgb <= "000000";
when "000111110001100" => rgb <= "000000";
when "000111110001101" => rgb <= "000000";
when "000111110001110" => rgb <= "000000";
when "000111110001111" => rgb <= "000000";
when "000111110010000" => rgb <= "000000";
when "000111110010001" => rgb <= "000000";
when "001000000001110" => rgb <= "000000";
when "001000000001111" => rgb <= "100110";
when "001000000010000" => rgb <= "100110";
when "001000000010001" => rgb <= "100110";
when "001000000010010" => rgb <= "100110";
when "001000000010011" => rgb <= "000000";
when "001000000010100" => rgb <= "000000";
when "001000000010101" => rgb <= "000000";
when "001000000010110" => rgb <= "000000";
when "001000000010111" => rgb <= "000000";
when "001000000011000" => rgb <= "000000";
when "001000000011001" => rgb <= "000000";
when "001000000011010" => rgb <= "000000";
when "001000000011011" => rgb <= "000000";
when "001000000011100" => rgb <= "000000";
when "001000000011101" => rgb <= "000000";
when "001000000011110" => rgb <= "000000";
when "001000000011111" => rgb <= "000000";
when "001000000100000" => rgb <= "000000";
when "001000000100001" => rgb <= "100110";
when "001000000100010" => rgb <= "100110";
when "001000000100011" => rgb <= "100110";
when "001000000100100" => rgb <= "000000";
when "001000000100101" => rgb <= "000000";
when "001000000100110" => rgb <= "000000";
when "001000000100111" => rgb <= "000000";
when "001000000101000" => rgb <= "000000";
when "001000000101001" => rgb <= "000000";
when "001000000101010" => rgb <= "100110";
when "001000000101011" => rgb <= "100110";
when "001000000101100" => rgb <= "100110";
when "001000000101101" => rgb <= "000000";
when "001000000101110" => rgb <= "000000";
when "001000000101111" => rgb <= "000000";
when "001000000110000" => rgb <= "000000";
when "001000000110001" => rgb <= "000000";
when "001000000110010" => rgb <= "000000";
when "001000000110011" => rgb <= "100110";
when "001000000110100" => rgb <= "100110";
when "001000000110101" => rgb <= "100110";
when "001000000110110" => rgb <= "000000";
when "001000000110111" => rgb <= "000000";
when "001000000111000" => rgb <= "100110";
when "001000000111001" => rgb <= "100110";
when "001000000111010" => rgb <= "100110";
when "001000000111011" => rgb <= "000000";
when "001000000111100" => rgb <= "000000";
when "001000000111101" => rgb <= "000000";
when "001000000111110" => rgb <= "000000";
when "001000000111111" => rgb <= "000000";
when "001000001000000" => rgb <= "100110";
when "001000001000001" => rgb <= "100110";
when "001000001000010" => rgb <= "100110";
when "001000001000011" => rgb <= "000000";
when "001000001000100" => rgb <= "000000";
when "001000001000101" => rgb <= "000000";
when "001000001000110" => rgb <= "000000";
when "001000001000111" => rgb <= "000000";
when "001000001001000" => rgb <= "000000";
when "001000001001001" => rgb <= "100110";
when "001000001001010" => rgb <= "100110";
when "001000001001011" => rgb <= "100110";
when "001000001001100" => rgb <= "000000";
when "001000001001101" => rgb <= "000000";
when "001000001001110" => rgb <= "000000";
when "001000001001111" => rgb <= "000000";
when "001000001010000" => rgb <= "000000";
when "001000001010001" => rgb <= "000000";
when "001000001010010" => rgb <= "000000";
when "001000001011001" => rgb <= "000000";
when "001000001011010" => rgb <= "100110";
when "001000001011011" => rgb <= "100110";
when "001000001011100" => rgb <= "100110";
when "001000001011101" => rgb <= "000000";
when "001000001011110" => rgb <= "000000";
when "001000001011111" => rgb <= "000000";
when "001000001100000" => rgb <= "000000";
when "001000001100001" => rgb <= "000000";
when "001000001100010" => rgb <= "000000";
when "001000001100011" => rgb <= "000000";
when "001000001100100" => rgb <= "000000";
when "001000001100101" => rgb <= "000000";
when "001000001100110" => rgb <= "000000";
when "001000001100111" => rgb <= "000000";
when "001000001101000" => rgb <= "100110";
when "001000001101001" => rgb <= "100110";
when "001000001101010" => rgb <= "100110";
when "001000001101011" => rgb <= "000000";
when "001000001101100" => rgb <= "000000";
when "001000001101101" => rgb <= "000000";
when "001000001101110" => rgb <= "000000";
when "001000001101111" => rgb <= "000000";
when "001000001110000" => rgb <= "000000";
when "001000001110001" => rgb <= "100110";
when "001000001110010" => rgb <= "100110";
when "001000001110011" => rgb <= "100110";
when "001000001110100" => rgb <= "000000";
when "001000001110101" => rgb <= "000000";
when "001000001110110" => rgb <= "100110";
when "001000001110111" => rgb <= "100110";
when "001000001111000" => rgb <= "100110";
when "001000001111001" => rgb <= "100110";
when "001000001111010" => rgb <= "100110";
when "001000001111011" => rgb <= "100110";
when "001000001111100" => rgb <= "100110";
when "001000001111101" => rgb <= "100110";
when "001000001111110" => rgb <= "100110";
when "001000001111111" => rgb <= "100110";
when "001000010000000" => rgb <= "100110";
when "001000010000001" => rgb <= "100110";
when "001000010000010" => rgb <= "100110";
when "001000010000011" => rgb <= "000000";
when "001000010000100" => rgb <= "000000";
when "001000010000101" => rgb <= "100110";
when "001000010000110" => rgb <= "100110";
when "001000010000111" => rgb <= "100110";
when "001000010001000" => rgb <= "000000";
when "001000010001001" => rgb <= "000000";
when "001000010001010" => rgb <= "000000";
when "001000010001011" => rgb <= "000000";
when "001000010001100" => rgb <= "000000";
when "001000010001101" => rgb <= "000000";
when "001000010001110" => rgb <= "000000";
when "001000010001111" => rgb <= "000000";
when "001000100001110" => rgb <= "000000";
when "001000100001111" => rgb <= "000000";
when "001000100010000" => rgb <= "000000";
when "001000100010001" => rgb <= "100110";
when "001000100010010" => rgb <= "100110";
when "001000100010011" => rgb <= "100110";
when "001000100010100" => rgb <= "100110";
when "001000100010101" => rgb <= "100110";
when "001000100010110" => rgb <= "100110";
when "001000100010111" => rgb <= "100110";
when "001000100011000" => rgb <= "100110";
when "001000100011001" => rgb <= "000000";
when "001000100011010" => rgb <= "000000";
when "001000100011011" => rgb <= "000000";
when "001000100011100" => rgb <= "000000";
when "001000100011101" => rgb <= "000000";
when "001000100100000" => rgb <= "000000";
when "001000100100001" => rgb <= "100110";
when "001000100100010" => rgb <= "100110";
when "001000100100011" => rgb <= "100110";
when "001000100100100" => rgb <= "000000";
when "001000100100101" => rgb <= "000000";
when "001000100100110" => rgb <= "000000";
when "001000100101001" => rgb <= "000000";
when "001000100101010" => rgb <= "100110";
when "001000100101011" => rgb <= "100110";
when "001000100101100" => rgb <= "100110";
when "001000100101101" => rgb <= "000000";
when "001000100101110" => rgb <= "000000";
when "001000100101111" => rgb <= "000000";
when "001000100110000" => rgb <= "000000";
when "001000100110001" => rgb <= "000000";
when "001000100110010" => rgb <= "000000";
when "001000100110011" => rgb <= "100110";
when "001000100110100" => rgb <= "100110";
when "001000100110101" => rgb <= "100110";
when "001000100110110" => rgb <= "000000";
when "001000100110111" => rgb <= "000000";
when "001000100111000" => rgb <= "100110";
when "001000100111001" => rgb <= "100110";
when "001000100111010" => rgb <= "100110";
when "001000100111011" => rgb <= "000000";
when "001000100111100" => rgb <= "000000";
when "001000100111101" => rgb <= "000000";
when "001000100111110" => rgb <= "000000";
when "001000100111111" => rgb <= "100110";
when "001000101000000" => rgb <= "100110";
when "001000101000001" => rgb <= "100110";
when "001000101000010" => rgb <= "100110";
when "001000101000011" => rgb <= "000000";
when "001000101000100" => rgb <= "000000";
when "001000101000101" => rgb <= "000000";
when "001000101001000" => rgb <= "000000";
when "001000101001001" => rgb <= "100110";
when "001000101001010" => rgb <= "100110";
when "001000101001011" => rgb <= "100110";
when "001000101001100" => rgb <= "000000";
when "001000101001101" => rgb <= "000000";
when "001000101001110" => rgb <= "000000";
when "001000101011001" => rgb <= "000000";
when "001000101011010" => rgb <= "100110";
when "001000101011011" => rgb <= "100110";
when "001000101011100" => rgb <= "100110";
when "001000101011101" => rgb <= "000000";
when "001000101011110" => rgb <= "000000";
when "001000101011111" => rgb <= "000000";
when "001000101100000" => rgb <= "100110";
when "001000101100001" => rgb <= "100110";
when "001000101100010" => rgb <= "100110";
when "001000101100011" => rgb <= "100110";
when "001000101100100" => rgb <= "100110";
when "001000101100101" => rgb <= "100110";
when "001000101100110" => rgb <= "000000";
when "001000101100111" => rgb <= "000000";
when "001000101101000" => rgb <= "100110";
when "001000101101001" => rgb <= "100110";
when "001000101101010" => rgb <= "100110";
when "001000101101011" => rgb <= "000000";
when "001000101101100" => rgb <= "000000";
when "001000101101101" => rgb <= "000000";
when "001000101101110" => rgb <= "000000";
when "001000101101111" => rgb <= "000000";
when "001000101110000" => rgb <= "000000";
when "001000101110001" => rgb <= "100110";
when "001000101110010" => rgb <= "100110";
when "001000101110011" => rgb <= "100110";
when "001000101110100" => rgb <= "000000";
when "001000101110101" => rgb <= "000000";
when "001000101110110" => rgb <= "100110";
when "001000101110111" => rgb <= "100110";
when "001000101111000" => rgb <= "100110";
when "001000101111001" => rgb <= "000000";
when "001000101111010" => rgb <= "100110";
when "001000101111011" => rgb <= "100110";
when "001000101111100" => rgb <= "100110";
when "001000101111101" => rgb <= "100110";
when "001000101111110" => rgb <= "100110";
when "001000101111111" => rgb <= "000000";
when "001000110000000" => rgb <= "100110";
when "001000110000001" => rgb <= "100110";
when "001000110000010" => rgb <= "100110";
when "001000110000011" => rgb <= "000000";
when "001000110000100" => rgb <= "000000";
when "001000110000101" => rgb <= "100110";
when "001000110000110" => rgb <= "100110";
when "001000110000111" => rgb <= "100110";
when "001000110001000" => rgb <= "100110";
when "001000110001001" => rgb <= "100110";
when "001000110001010" => rgb <= "100110";
when "001000110001011" => rgb <= "100110";
when "001000110001100" => rgb <= "100110";
when "001000110001101" => rgb <= "100110";
when "001000110001110" => rgb <= "000000";
when "001000110001111" => rgb <= "000000";
when "001001000010000" => rgb <= "000000";
when "001001000010001" => rgb <= "100110";
when "001001000010010" => rgb <= "100110";
when "001001000010011" => rgb <= "100110";
when "001001000010100" => rgb <= "100110";
when "001001000010101" => rgb <= "100110";
when "001001000010110" => rgb <= "100110";
when "001001000010111" => rgb <= "100110";
when "001001000011000" => rgb <= "100110";
when "001001000011001" => rgb <= "100110";
when "001001000011010" => rgb <= "100110";
when "001001000011011" => rgb <= "000000";
when "001001000011100" => rgb <= "000000";
when "001001000011101" => rgb <= "000000";
when "001001000100000" => rgb <= "000000";
when "001001000100001" => rgb <= "100110";
when "001001000100010" => rgb <= "100110";
when "001001000100011" => rgb <= "100110";
when "001001000100100" => rgb <= "000000";
when "001001000100101" => rgb <= "000000";
when "001001000100110" => rgb <= "000000";
when "001001000101001" => rgb <= "000000";
when "001001000101010" => rgb <= "100110";
when "001001000101011" => rgb <= "100110";
when "001001000101100" => rgb <= "100110";
when "001001000101101" => rgb <= "100110";
when "001001000101110" => rgb <= "100110";
when "001001000101111" => rgb <= "100110";
when "001001000110000" => rgb <= "100110";
when "001001000110001" => rgb <= "100110";
when "001001000110010" => rgb <= "100110";
when "001001000110011" => rgb <= "100110";
when "001001000110100" => rgb <= "100110";
when "001001000110101" => rgb <= "100110";
when "001001000110110" => rgb <= "000000";
when "001001000110111" => rgb <= "000000";
when "001001000111000" => rgb <= "100110";
when "001001000111001" => rgb <= "100110";
when "001001000111010" => rgb <= "100110";
when "001001000111011" => rgb <= "100110";
when "001001000111100" => rgb <= "100110";
when "001001000111101" => rgb <= "100110";
when "001001000111110" => rgb <= "100110";
when "001001000111111" => rgb <= "100110";
when "001001001000000" => rgb <= "100110";
when "001001001000001" => rgb <= "000000";
when "001001001000010" => rgb <= "000000";
when "001001001000011" => rgb <= "000000";
when "001001001000100" => rgb <= "000000";
when "001001001001000" => rgb <= "000000";
when "001001001001001" => rgb <= "100110";
when "001001001001010" => rgb <= "100110";
when "001001001001011" => rgb <= "100110";
when "001001001001100" => rgb <= "000000";
when "001001001001101" => rgb <= "000000";
when "001001001001110" => rgb <= "000000";
when "001001001011001" => rgb <= "000000";
when "001001001011010" => rgb <= "100110";
when "001001001011011" => rgb <= "100110";
when "001001001011100" => rgb <= "100110";
when "001001001011101" => rgb <= "000000";
when "001001001011110" => rgb <= "000000";
when "001001001011111" => rgb <= "000000";
when "001001001100000" => rgb <= "100110";
when "001001001100001" => rgb <= "100110";
when "001001001100010" => rgb <= "100110";
when "001001001100011" => rgb <= "100110";
when "001001001100100" => rgb <= "100110";
when "001001001100101" => rgb <= "100110";
when "001001001100110" => rgb <= "000000";
when "001001001100111" => rgb <= "000000";
when "001001001101000" => rgb <= "100110";
when "001001001101001" => rgb <= "100110";
when "001001001101010" => rgb <= "100110";
when "001001001101011" => rgb <= "100110";
when "001001001101100" => rgb <= "100110";
when "001001001101101" => rgb <= "100110";
when "001001001101110" => rgb <= "100110";
when "001001001101111" => rgb <= "100110";
when "001001001110000" => rgb <= "100110";
when "001001001110001" => rgb <= "100110";
when "001001001110010" => rgb <= "100110";
when "001001001110011" => rgb <= "100110";
when "001001001110100" => rgb <= "000000";
when "001001001110101" => rgb <= "000000";
when "001001001110110" => rgb <= "100110";
when "001001001110111" => rgb <= "100110";
when "001001001111000" => rgb <= "100110";
when "001001001111001" => rgb <= "000000";
when "001001001111010" => rgb <= "100110";
when "001001001111011" => rgb <= "100110";
when "001001001111100" => rgb <= "100110";
when "001001001111101" => rgb <= "100110";
when "001001001111110" => rgb <= "100110";
when "001001001111111" => rgb <= "000000";
when "001001010000000" => rgb <= "100110";
when "001001010000001" => rgb <= "100110";
when "001001010000010" => rgb <= "100110";
when "001001010000011" => rgb <= "000000";
when "001001010000100" => rgb <= "000000";
when "001001010000101" => rgb <= "100110";
when "001001010000110" => rgb <= "100110";
when "001001010000111" => rgb <= "100110";
when "001001010001000" => rgb <= "100110";
when "001001010001001" => rgb <= "100110";
when "001001010001010" => rgb <= "100110";
when "001001010001011" => rgb <= "100110";
when "001001010001100" => rgb <= "100110";
when "001001010001101" => rgb <= "100110";
when "001001010001110" => rgb <= "000000";
when "001001010001111" => rgb <= "000000";
when "001001100001110" => rgb <= "000000";
when "001001100001111" => rgb <= "000000";
when "001001100010000" => rgb <= "000000";
when "001001100010001" => rgb <= "000000";
when "001001100010010" => rgb <= "000000";
when "001001100010011" => rgb <= "000000";
when "001001100010100" => rgb <= "000000";
when "001001100010101" => rgb <= "000000";
when "001001100010110" => rgb <= "000000";
when "001001100010111" => rgb <= "100110";
when "001001100011000" => rgb <= "100110";
when "001001100011001" => rgb <= "100110";
when "001001100011010" => rgb <= "100110";
when "001001100011011" => rgb <= "000000";
when "001001100011100" => rgb <= "000000";
when "001001100011101" => rgb <= "000000";
when "001001100100000" => rgb <= "000000";
when "001001100100001" => rgb <= "100110";
when "001001100100010" => rgb <= "100110";
when "001001100100011" => rgb <= "100110";
when "001001100100100" => rgb <= "000000";
when "001001100100101" => rgb <= "000000";
when "001001100100110" => rgb <= "000000";
when "001001100101001" => rgb <= "000000";
when "001001100101010" => rgb <= "100110";
when "001001100101011" => rgb <= "100110";
when "001001100101100" => rgb <= "100110";
when "001001100101101" => rgb <= "100110";
when "001001100101110" => rgb <= "100110";
when "001001100101111" => rgb <= "100110";
when "001001100110000" => rgb <= "100110";
when "001001100110001" => rgb <= "100110";
when "001001100110010" => rgb <= "100110";
when "001001100110011" => rgb <= "100110";
when "001001100110100" => rgb <= "100110";
when "001001100110101" => rgb <= "100110";
when "001001100110110" => rgb <= "000000";
when "001001100110111" => rgb <= "000000";
when "001001100111000" => rgb <= "100110";
when "001001100111001" => rgb <= "100110";
when "001001100111010" => rgb <= "100110";
when "001001100111011" => rgb <= "100110";
when "001001100111100" => rgb <= "100110";
when "001001100111101" => rgb <= "100110";
when "001001100111110" => rgb <= "100110";
when "001001100111111" => rgb <= "100110";
when "001001101000000" => rgb <= "000000";
when "001001101000001" => rgb <= "000000";
when "001001101000010" => rgb <= "000000";
when "001001101000011" => rgb <= "000000";
when "001001101001000" => rgb <= "000000";
when "001001101001001" => rgb <= "100110";
when "001001101001010" => rgb <= "100110";
when "001001101001011" => rgb <= "100110";
when "001001101001100" => rgb <= "000000";
when "001001101001101" => rgb <= "000000";
when "001001101001110" => rgb <= "000000";
when "001001101011001" => rgb <= "000000";
when "001001101011010" => rgb <= "100110";
when "001001101011011" => rgb <= "100110";
when "001001101011100" => rgb <= "100110";
when "001001101011101" => rgb <= "000000";
when "001001101011110" => rgb <= "000000";
when "001001101011111" => rgb <= "000000";
when "001001101100000" => rgb <= "000000";
when "001001101100001" => rgb <= "000000";
when "001001101100010" => rgb <= "000000";
when "001001101100011" => rgb <= "100110";
when "001001101100100" => rgb <= "100110";
when "001001101100101" => rgb <= "100110";
when "001001101100110" => rgb <= "000000";
when "001001101100111" => rgb <= "000000";
when "001001101101000" => rgb <= "100110";
when "001001101101001" => rgb <= "100110";
when "001001101101010" => rgb <= "100110";
when "001001101101011" => rgb <= "100110";
when "001001101101100" => rgb <= "100110";
when "001001101101101" => rgb <= "100110";
when "001001101101110" => rgb <= "100110";
when "001001101101111" => rgb <= "100110";
when "001001101110000" => rgb <= "100110";
when "001001101110001" => rgb <= "100110";
when "001001101110010" => rgb <= "100110";
when "001001101110011" => rgb <= "100110";
when "001001101110100" => rgb <= "000000";
when "001001101110101" => rgb <= "000000";
when "001001101110110" => rgb <= "100110";
when "001001101110111" => rgb <= "100110";
when "001001101111000" => rgb <= "100110";
when "001001101111001" => rgb <= "000000";
when "001001101111010" => rgb <= "000000";
when "001001101111011" => rgb <= "100110";
when "001001101111100" => rgb <= "100110";
when "001001101111101" => rgb <= "100110";
when "001001101111110" => rgb <= "000000";
when "001001101111111" => rgb <= "000000";
when "001001110000000" => rgb <= "100110";
when "001001110000001" => rgb <= "100110";
when "001001110000010" => rgb <= "100110";
when "001001110000011" => rgb <= "000000";
when "001001110000100" => rgb <= "000000";
when "001001110000101" => rgb <= "100110";
when "001001110000110" => rgb <= "100110";
when "001001110000111" => rgb <= "100110";
when "001001110001000" => rgb <= "000000";
when "001001110001001" => rgb <= "000000";
when "001001110001010" => rgb <= "000000";
when "001001110001011" => rgb <= "000000";
when "001001110001100" => rgb <= "000000";
when "001001110001101" => rgb <= "000000";
when "001001110001110" => rgb <= "000000";
when "001001110001111" => rgb <= "000000";
when "001010000001110" => rgb <= "000000";
when "001010000001111" => rgb <= "100110";
when "001010000010000" => rgb <= "100110";
when "001010000010001" => rgb <= "100110";
when "001010000010010" => rgb <= "100110";
when "001010000010011" => rgb <= "000000";
when "001010000010100" => rgb <= "000000";
when "001010000010101" => rgb <= "000000";
when "001010000010110" => rgb <= "000000";
when "001010000010111" => rgb <= "100110";
when "001010000011000" => rgb <= "100110";
when "001010000011001" => rgb <= "100110";
when "001010000011010" => rgb <= "100110";
when "001010000011011" => rgb <= "000000";
when "001010000011100" => rgb <= "000000";
when "001010000011101" => rgb <= "000000";
when "001010000100000" => rgb <= "000000";
when "001010000100001" => rgb <= "100110";
when "001010000100010" => rgb <= "100110";
when "001010000100011" => rgb <= "100110";
when "001010000100100" => rgb <= "000000";
when "001010000100101" => rgb <= "000000";
when "001010000100110" => rgb <= "000000";
when "001010000101001" => rgb <= "000000";
when "001010000101010" => rgb <= "100110";
when "001010000101011" => rgb <= "100110";
when "001010000101100" => rgb <= "100110";
when "001010000101101" => rgb <= "000000";
when "001010000101110" => rgb <= "000000";
when "001010000101111" => rgb <= "000000";
when "001010000110000" => rgb <= "000000";
when "001010000110001" => rgb <= "000000";
when "001010000110010" => rgb <= "000000";
when "001010000110011" => rgb <= "100110";
when "001010000110100" => rgb <= "100110";
when "001010000110101" => rgb <= "100110";
when "001010000110110" => rgb <= "000000";
when "001010000110111" => rgb <= "000000";
when "001010000111000" => rgb <= "100110";
when "001010000111001" => rgb <= "100110";
when "001010000111010" => rgb <= "100110";
when "001010000111011" => rgb <= "000000";
when "001010000111100" => rgb <= "000000";
when "001010000111101" => rgb <= "100110";
when "001010000111110" => rgb <= "100110";
when "001010000111111" => rgb <= "100110";
when "001010001000000" => rgb <= "100110";
when "001010001000001" => rgb <= "000000";
when "001010001000010" => rgb <= "000000";
when "001010001000011" => rgb <= "000000";
when "001010001000100" => rgb <= "000000";
when "001010001001000" => rgb <= "000000";
when "001010001001001" => rgb <= "100110";
when "001010001001010" => rgb <= "100110";
when "001010001001011" => rgb <= "100110";
when "001010001001100" => rgb <= "000000";
when "001010001001101" => rgb <= "000000";
when "001010001001110" => rgb <= "000000";
when "001010001011001" => rgb <= "000000";
when "001010001011010" => rgb <= "100110";
when "001010001011011" => rgb <= "100110";
when "001010001011100" => rgb <= "100110";
when "001010001011101" => rgb <= "000000";
when "001010001011110" => rgb <= "000000";
when "001010001011111" => rgb <= "000000";
when "001010001100000" => rgb <= "000000";
when "001010001100001" => rgb <= "000000";
when "001010001100010" => rgb <= "000000";
when "001010001100011" => rgb <= "100110";
when "001010001100100" => rgb <= "100110";
when "001010001100101" => rgb <= "100110";
when "001010001100110" => rgb <= "000000";
when "001010001100111" => rgb <= "000000";
when "001010001101000" => rgb <= "100110";
when "001010001101001" => rgb <= "100110";
when "001010001101010" => rgb <= "100110";
when "001010001101011" => rgb <= "000000";
when "001010001101100" => rgb <= "000000";
when "001010001101101" => rgb <= "000000";
when "001010001101110" => rgb <= "000000";
when "001010001101111" => rgb <= "000000";
when "001010001110000" => rgb <= "000000";
when "001010001110001" => rgb <= "100110";
when "001010001110010" => rgb <= "100110";
when "001010001110011" => rgb <= "100110";
when "001010001110100" => rgb <= "000000";
when "001010001110101" => rgb <= "000000";
when "001010001110110" => rgb <= "100110";
when "001010001110111" => rgb <= "100110";
when "001010001111000" => rgb <= "100110";
when "001010001111001" => rgb <= "000000";
when "001010001111010" => rgb <= "000000";
when "001010001111011" => rgb <= "100110";
when "001010001111100" => rgb <= "100110";
when "001010001111101" => rgb <= "100110";
when "001010001111110" => rgb <= "000000";
when "001010001111111" => rgb <= "000000";
when "001010010000000" => rgb <= "100110";
when "001010010000001" => rgb <= "100110";
when "001010010000010" => rgb <= "100110";
when "001010010000011" => rgb <= "000000";
when "001010010000100" => rgb <= "000000";
when "001010010000101" => rgb <= "100110";
when "001010010000110" => rgb <= "100110";
when "001010010000111" => rgb <= "100110";
when "001010010001000" => rgb <= "000000";
when "001010010001001" => rgb <= "000000";
when "001010010001010" => rgb <= "000000";
when "001010010001011" => rgb <= "000000";
when "001010010001100" => rgb <= "000000";
when "001010010001101" => rgb <= "000000";
when "001010010001110" => rgb <= "000000";
when "001010010001111" => rgb <= "000000";
when "001010100001110" => rgb <= "000000";
when "001010100001111" => rgb <= "100110";
when "001010100010000" => rgb <= "100110";
when "001010100010001" => rgb <= "100110";
when "001010100010010" => rgb <= "100110";
when "001010100010011" => rgb <= "000000";
when "001010100010100" => rgb <= "000000";
when "001010100010101" => rgb <= "000000";
when "001010100010110" => rgb <= "000000";
when "001010100010111" => rgb <= "100110";
when "001010100011000" => rgb <= "100110";
when "001010100011001" => rgb <= "100110";
when "001010100011010" => rgb <= "100110";
when "001010100011011" => rgb <= "000000";
when "001010100011100" => rgb <= "000000";
when "001010100011101" => rgb <= "000000";
when "001010100100000" => rgb <= "000000";
when "001010100100001" => rgb <= "100110";
when "001010100100010" => rgb <= "100110";
when "001010100100011" => rgb <= "100110";
when "001010100100100" => rgb <= "000000";
when "001010100100101" => rgb <= "000000";
when "001010100100110" => rgb <= "000000";
when "001010100101001" => rgb <= "000000";
when "001010100101010" => rgb <= "100110";
when "001010100101011" => rgb <= "100110";
when "001010100101100" => rgb <= "100110";
when "001010100101101" => rgb <= "000000";
when "001010100101110" => rgb <= "000000";
when "001010100101111" => rgb <= "000000";
when "001010100110000" => rgb <= "000000";
when "001010100110001" => rgb <= "000000";
when "001010100110010" => rgb <= "000000";
when "001010100110011" => rgb <= "100110";
when "001010100110100" => rgb <= "100110";
when "001010100110101" => rgb <= "100110";
when "001010100110110" => rgb <= "000000";
when "001010100110111" => rgb <= "000000";
when "001010100111000" => rgb <= "100110";
when "001010100111001" => rgb <= "100110";
when "001010100111010" => rgb <= "100110";
when "001010100111011" => rgb <= "000000";
when "001010100111100" => rgb <= "000000";
when "001010100111101" => rgb <= "000000";
when "001010100111110" => rgb <= "100110";
when "001010100111111" => rgb <= "100110";
when "001010101000000" => rgb <= "100110";
when "001010101000001" => rgb <= "100110";
when "001010101000010" => rgb <= "000000";
when "001010101000011" => rgb <= "000000";
when "001010101000100" => rgb <= "000000";
when "001010101001000" => rgb <= "000000";
when "001010101001001" => rgb <= "100110";
when "001010101001010" => rgb <= "100110";
when "001010101001011" => rgb <= "100110";
when "001010101001100" => rgb <= "000000";
when "001010101001101" => rgb <= "000000";
when "001010101001110" => rgb <= "000000";
when "001010101011001" => rgb <= "000000";
when "001010101011010" => rgb <= "100110";
when "001010101011011" => rgb <= "100110";
when "001010101011100" => rgb <= "100110";
when "001010101011101" => rgb <= "100110";
when "001010101011110" => rgb <= "000000";
when "001010101011111" => rgb <= "000000";
when "001010101100000" => rgb <= "000000";
when "001010101100001" => rgb <= "000000";
when "001010101100010" => rgb <= "000000";
when "001010101100011" => rgb <= "100110";
when "001010101100100" => rgb <= "100110";
when "001010101100101" => rgb <= "100110";
when "001010101100110" => rgb <= "000000";
when "001010101100111" => rgb <= "000000";
when "001010101101000" => rgb <= "100110";
when "001010101101001" => rgb <= "100110";
when "001010101101010" => rgb <= "100110";
when "001010101101011" => rgb <= "000000";
when "001010101101100" => rgb <= "000000";
when "001010101101101" => rgb <= "000000";
when "001010101101110" => rgb <= "000000";
when "001010101101111" => rgb <= "000000";
when "001010101110000" => rgb <= "000000";
when "001010101110001" => rgb <= "100110";
when "001010101110010" => rgb <= "100110";
when "001010101110011" => rgb <= "100110";
when "001010101110100" => rgb <= "000000";
when "001010101110101" => rgb <= "000000";
when "001010101110110" => rgb <= "100110";
when "001010101110111" => rgb <= "100110";
when "001010101111000" => rgb <= "100110";
when "001010101111001" => rgb <= "000000";
when "001010101111010" => rgb <= "000000";
when "001010101111011" => rgb <= "100110";
when "001010101111100" => rgb <= "100110";
when "001010101111101" => rgb <= "100110";
when "001010101111110" => rgb <= "000000";
when "001010101111111" => rgb <= "000000";
when "001010110000000" => rgb <= "100110";
when "001010110000001" => rgb <= "100110";
when "001010110000010" => rgb <= "100110";
when "001010110000011" => rgb <= "000000";
when "001010110000100" => rgb <= "000000";
when "001010110000101" => rgb <= "100110";
when "001010110000110" => rgb <= "100110";
when "001010110000111" => rgb <= "100110";
when "001010110001000" => rgb <= "000000";
when "001010110001001" => rgb <= "000000";
when "001010110001010" => rgb <= "000000";
when "001010110001011" => rgb <= "000000";
when "001010110001100" => rgb <= "000000";
when "001010110001101" => rgb <= "000000";
when "001010110001110" => rgb <= "000000";
when "001010110001111" => rgb <= "000000";
when "001011000001110" => rgb <= "000000";
when "001011000001111" => rgb <= "100110";
when "001011000010000" => rgb <= "100110";
when "001011000010001" => rgb <= "100110";
when "001011000010010" => rgb <= "100110";
when "001011000010011" => rgb <= "100110";
when "001011000010100" => rgb <= "100110";
when "001011000010101" => rgb <= "100110";
when "001011000010110" => rgb <= "100110";
when "001011000010111" => rgb <= "100110";
when "001011000011000" => rgb <= "100110";
when "001011000011001" => rgb <= "100110";
when "001011000011010" => rgb <= "100110";
when "001011000011011" => rgb <= "000000";
when "001011000011100" => rgb <= "000000";
when "001011000011101" => rgb <= "000000";
when "001011000100000" => rgb <= "000000";
when "001011000100001" => rgb <= "100110";
when "001011000100010" => rgb <= "100110";
when "001011000100011" => rgb <= "100110";
when "001011000100100" => rgb <= "000000";
when "001011000100101" => rgb <= "000000";
when "001011000100110" => rgb <= "000000";
when "001011000101001" => rgb <= "000000";
when "001011000101010" => rgb <= "100110";
when "001011000101011" => rgb <= "100110";
when "001011000101100" => rgb <= "100110";
when "001011000101101" => rgb <= "000000";
when "001011000101110" => rgb <= "000000";
when "001011000101111" => rgb <= "000000";
when "001011000110000" => rgb <= "000000";
when "001011000110001" => rgb <= "000000";
when "001011000110010" => rgb <= "000000";
when "001011000110011" => rgb <= "100110";
when "001011000110100" => rgb <= "100110";
when "001011000110101" => rgb <= "100110";
when "001011000110110" => rgb <= "000000";
when "001011000110111" => rgb <= "000000";
when "001011000111000" => rgb <= "100110";
when "001011000111001" => rgb <= "100110";
when "001011000111010" => rgb <= "100110";
when "001011000111011" => rgb <= "000000";
when "001011000111100" => rgb <= "000000";
when "001011000111101" => rgb <= "000000";
when "001011000111110" => rgb <= "000000";
when "001011000111111" => rgb <= "100110";
when "001011001000000" => rgb <= "100110";
when "001011001000001" => rgb <= "100110";
when "001011001000010" => rgb <= "000000";
when "001011001000011" => rgb <= "000000";
when "001011001000100" => rgb <= "000000";
when "001011001001000" => rgb <= "000000";
when "001011001001001" => rgb <= "100110";
when "001011001001010" => rgb <= "100110";
when "001011001001011" => rgb <= "100110";
when "001011001001100" => rgb <= "000000";
when "001011001001101" => rgb <= "000000";
when "001011001001110" => rgb <= "000000";
when "001011001011001" => rgb <= "000000";
when "001011001011010" => rgb <= "100110";
when "001011001011011" => rgb <= "100110";
when "001011001011100" => rgb <= "100110";
when "001011001011101" => rgb <= "100110";
when "001011001011110" => rgb <= "100110";
when "001011001011111" => rgb <= "100110";
when "001011001100000" => rgb <= "100110";
when "001011001100001" => rgb <= "100110";
when "001011001100010" => rgb <= "100110";
when "001011001100011" => rgb <= "100110";
when "001011001100100" => rgb <= "100110";
when "001011001100101" => rgb <= "100110";
when "001011001100110" => rgb <= "000000";
when "001011001100111" => rgb <= "000000";
when "001011001101000" => rgb <= "100110";
when "001011001101001" => rgb <= "100110";
when "001011001101010" => rgb <= "100110";
when "001011001101011" => rgb <= "000000";
when "001011001101100" => rgb <= "000000";
when "001011001101101" => rgb <= "000000";
when "001011001101110" => rgb <= "000000";
when "001011001101111" => rgb <= "000000";
when "001011001110000" => rgb <= "000000";
when "001011001110001" => rgb <= "100110";
when "001011001110010" => rgb <= "100110";
when "001011001110011" => rgb <= "100110";
when "001011001110100" => rgb <= "000000";
when "001011001110101" => rgb <= "000000";
when "001011001110110" => rgb <= "100110";
when "001011001110111" => rgb <= "100110";
when "001011001111000" => rgb <= "100110";
when "001011001111001" => rgb <= "000000";
when "001011001111010" => rgb <= "000000";
when "001011001111011" => rgb <= "000000";
when "001011001111100" => rgb <= "000000";
when "001011001111101" => rgb <= "000000";
when "001011001111110" => rgb <= "000000";
when "001011001111111" => rgb <= "000000";
when "001011010000000" => rgb <= "100110";
when "001011010000001" => rgb <= "100110";
when "001011010000010" => rgb <= "100110";
when "001011010000011" => rgb <= "000000";
when "001011010000100" => rgb <= "000000";
when "001011010000101" => rgb <= "100110";
when "001011010000110" => rgb <= "100110";
when "001011010000111" => rgb <= "100110";
when "001011010001000" => rgb <= "100110";
when "001011010001001" => rgb <= "100110";
when "001011010001010" => rgb <= "100110";
when "001011010001011" => rgb <= "100110";
when "001011010001100" => rgb <= "100110";
when "001011010001101" => rgb <= "100110";
when "001011010001110" => rgb <= "100110";
when "001011010001111" => rgb <= "000000";
when "001011010010000" => rgb <= "000000";
when "001011010010001" => rgb <= "000000";
when "001011100001110" => rgb <= "000000";
when "001011100001111" => rgb <= "000000";
when "001011100010000" => rgb <= "000000";
when "001011100010001" => rgb <= "100110";
when "001011100010010" => rgb <= "100110";
when "001011100010011" => rgb <= "100110";
when "001011100010100" => rgb <= "100110";
when "001011100010101" => rgb <= "100110";
when "001011100010110" => rgb <= "100110";
when "001011100010111" => rgb <= "100110";
when "001011100011000" => rgb <= "100110";
when "001011100011001" => rgb <= "000000";
when "001011100011010" => rgb <= "000000";
when "001011100011011" => rgb <= "000000";
when "001011100011100" => rgb <= "000000";
when "001011100011101" => rgb <= "000000";
when "001011100100000" => rgb <= "000000";
when "001011100100001" => rgb <= "100110";
when "001011100100010" => rgb <= "100110";
when "001011100100011" => rgb <= "100110";
when "001011100100100" => rgb <= "000000";
when "001011100100101" => rgb <= "000000";
when "001011100100110" => rgb <= "000000";
when "001011100101001" => rgb <= "000000";
when "001011100101010" => rgb <= "100110";
when "001011100101011" => rgb <= "100110";
when "001011100101100" => rgb <= "100110";
when "001011100101101" => rgb <= "000000";
when "001011100101110" => rgb <= "000000";
when "001011100101111" => rgb <= "000000";
when "001011100110010" => rgb <= "000000";
when "001011100110011" => rgb <= "100110";
when "001011100110100" => rgb <= "100110";
when "001011100110101" => rgb <= "100110";
when "001011100110110" => rgb <= "000000";
when "001011100110111" => rgb <= "000000";
when "001011100111000" => rgb <= "100110";
when "001011100111001" => rgb <= "100110";
when "001011100111010" => rgb <= "100110";
when "001011100111011" => rgb <= "000000";
when "001011100111100" => rgb <= "000000";
when "001011100111101" => rgb <= "000000";
when "001011100111110" => rgb <= "000000";
when "001011100111111" => rgb <= "100110";
when "001011101000000" => rgb <= "100110";
when "001011101000001" => rgb <= "100110";
when "001011101000010" => rgb <= "000000";
when "001011101000011" => rgb <= "000000";
when "001011101000100" => rgb <= "000000";
when "001011101001000" => rgb <= "000000";
when "001011101001001" => rgb <= "100110";
when "001011101001010" => rgb <= "100110";
when "001011101001011" => rgb <= "100110";
when "001011101001100" => rgb <= "000000";
when "001011101001101" => rgb <= "000000";
when "001011101001110" => rgb <= "000000";
when "001011101011001" => rgb <= "000000";
when "001011101011010" => rgb <= "000000";
when "001011101011011" => rgb <= "100110";
when "001011101011100" => rgb <= "100110";
when "001011101011101" => rgb <= "100110";
when "001011101011110" => rgb <= "100110";
when "001011101011111" => rgb <= "100110";
when "001011101100000" => rgb <= "100110";
when "001011101100001" => rgb <= "100110";
when "001011101100010" => rgb <= "100110";
when "001011101100011" => rgb <= "100110";
when "001011101100100" => rgb <= "100110";
when "001011101100101" => rgb <= "100110";
when "001011101100110" => rgb <= "000000";
when "001011101100111" => rgb <= "000000";
when "001011101101000" => rgb <= "100110";
when "001011101101001" => rgb <= "100110";
when "001011101101010" => rgb <= "100110";
when "001011101101011" => rgb <= "000000";
when "001011101101100" => rgb <= "000000";
when "001011101101101" => rgb <= "000000";
when "001011101110000" => rgb <= "000000";
when "001011101110001" => rgb <= "100110";
when "001011101110010" => rgb <= "100110";
when "001011101110011" => rgb <= "100110";
when "001011101110100" => rgb <= "000000";
when "001011101110101" => rgb <= "000000";
when "001011101110110" => rgb <= "100110";
when "001011101110111" => rgb <= "100110";
when "001011101111000" => rgb <= "100110";
when "001011101111001" => rgb <= "000000";
when "001011101111010" => rgb <= "000000";
when "001011101111011" => rgb <= "000000";
when "001011101111100" => rgb <= "000000";
when "001011101111101" => rgb <= "000000";
when "001011101111110" => rgb <= "000000";
when "001011101111111" => rgb <= "000000";
when "001011110000000" => rgb <= "100110";
when "001011110000001" => rgb <= "100110";
when "001011110000010" => rgb <= "100110";
when "001011110000011" => rgb <= "000000";
when "001011110000100" => rgb <= "000000";
when "001011110000101" => rgb <= "100110";
when "001011110000110" => rgb <= "100110";
when "001011110000111" => rgb <= "100110";
when "001011110001000" => rgb <= "100110";
when "001011110001001" => rgb <= "100110";
when "001011110001010" => rgb <= "100110";
when "001011110001011" => rgb <= "100110";
when "001011110001100" => rgb <= "100110";
when "001011110001101" => rgb <= "100110";
when "001011110001110" => rgb <= "100110";
when "001011110001111" => rgb <= "000000";
when "001011110010000" => rgb <= "000000";
when "001011110010001" => rgb <= "000000";
when "001100000001111" => rgb <= "000000";
when "001100000010000" => rgb <= "000000";
when "001100000010001" => rgb <= "100110";
when "001100000010010" => rgb <= "100110";
when "001100000010011" => rgb <= "100110";
when "001100000010100" => rgb <= "100110";
when "001100000010101" => rgb <= "100110";
when "001100000010110" => rgb <= "100110";
when "001100000010111" => rgb <= "100110";
when "001100000011000" => rgb <= "100110";
when "001100000011001" => rgb <= "000000";
when "001100000011010" => rgb <= "000000";
when "001100000011011" => rgb <= "000000";
when "001100000011100" => rgb <= "000000";
when "001100000100000" => rgb <= "000000";
when "001100000100001" => rgb <= "100110";
when "001100000100010" => rgb <= "100110";
when "001100000100011" => rgb <= "100110";
when "001100000100100" => rgb <= "000000";
when "001100000100101" => rgb <= "000000";
when "001100000100110" => rgb <= "000000";
when "001100000101001" => rgb <= "000000";
when "001100000101010" => rgb <= "100110";
when "001100000101011" => rgb <= "100110";
when "001100000101100" => rgb <= "100110";
when "001100000101101" => rgb <= "000000";
when "001100000101110" => rgb <= "000000";
when "001100000101111" => rgb <= "000000";
when "001100000110010" => rgb <= "000000";
when "001100000110011" => rgb <= "100110";
when "001100000110100" => rgb <= "100110";
when "001100000110101" => rgb <= "100110";
when "001100000110110" => rgb <= "000000";
when "001100000110111" => rgb <= "000000";
when "001100000111000" => rgb <= "100110";
when "001100000111001" => rgb <= "100110";
when "001100000111010" => rgb <= "100110";
when "001100000111011" => rgb <= "000000";
when "001100000111100" => rgb <= "000000";
when "001100000111101" => rgb <= "000000";
when "001100000111110" => rgb <= "000000";
when "001100000111111" => rgb <= "100110";
when "001100001000000" => rgb <= "100110";
when "001100001000001" => rgb <= "100110";
when "001100001000010" => rgb <= "000000";
when "001100001000011" => rgb <= "000000";
when "001100001000100" => rgb <= "000000";
when "001100001001000" => rgb <= "000000";
when "001100001001001" => rgb <= "100110";
when "001100001001010" => rgb <= "100110";
when "001100001001011" => rgb <= "100110";
when "001100001001100" => rgb <= "000000";
when "001100001001101" => rgb <= "000000";
when "001100001001110" => rgb <= "000000";
when "001100001011010" => rgb <= "000000";
when "001100001011011" => rgb <= "000000";
when "001100001011100" => rgb <= "000000";
when "001100001011101" => rgb <= "100110";
when "001100001011110" => rgb <= "100110";
when "001100001011111" => rgb <= "100110";
when "001100001100000" => rgb <= "100110";
when "001100001100001" => rgb <= "100110";
when "001100001100010" => rgb <= "100110";
when "001100001100011" => rgb <= "100110";
when "001100001100100" => rgb <= "100110";
when "001100001100101" => rgb <= "100110";
when "001100001100110" => rgb <= "000000";
when "001100001100111" => rgb <= "000000";
when "001100001101000" => rgb <= "100110";
when "001100001101001" => rgb <= "100110";
when "001100001101010" => rgb <= "100110";
when "001100001101011" => rgb <= "000000";
when "001100001101100" => rgb <= "000000";
when "001100001101101" => rgb <= "000000";
when "001100001110000" => rgb <= "000000";
when "001100001110001" => rgb <= "100110";
when "001100001110010" => rgb <= "100110";
when "001100001110011" => rgb <= "100110";
when "001100001110100" => rgb <= "000000";
when "001100001110101" => rgb <= "000000";
when "001100001110110" => rgb <= "100110";
when "001100001110111" => rgb <= "100110";
when "001100001111000" => rgb <= "100110";
when "001100001111001" => rgb <= "000000";
when "001100001111010" => rgb <= "000000";
when "001100001111100" => rgb <= "000000";
when "001100001111101" => rgb <= "000000";
when "001100001111110" => rgb <= "000000";
when "001100001111111" => rgb <= "000000";
when "001100010000000" => rgb <= "100110";
when "001100010000001" => rgb <= "100110";
when "001100010000010" => rgb <= "100110";
when "001100010000011" => rgb <= "000000";
when "001100010000100" => rgb <= "000000";
when "001100010000101" => rgb <= "100110";
when "001100010000110" => rgb <= "100110";
when "001100010000111" => rgb <= "100110";
when "001100010001000" => rgb <= "100110";
when "001100010001001" => rgb <= "100110";
when "001100010001010" => rgb <= "100110";
when "001100010001011" => rgb <= "100110";
when "001100010001100" => rgb <= "100110";
when "001100010001101" => rgb <= "100110";
when "001100010001110" => rgb <= "100110";
when "001100010001111" => rgb <= "000000";
when "001100010010000" => rgb <= "000000";
when "001100010010001" => rgb <= "000000";
when "001100100001111" => rgb <= "000000";
when "001100100010000" => rgb <= "000000";
when "001100100010001" => rgb <= "000000";
when "001100100010010" => rgb <= "000000";
when "001100100010011" => rgb <= "000000";
when "001100100010100" => rgb <= "000000";
when "001100100010101" => rgb <= "000000";
when "001100100010110" => rgb <= "000000";
when "001100100010111" => rgb <= "000000";
when "001100100011000" => rgb <= "000000";
when "001100100011001" => rgb <= "000000";
when "001100100011010" => rgb <= "000000";
when "001100100011011" => rgb <= "000000";
when "001100100011100" => rgb <= "000000";
when "001100100100000" => rgb <= "000000";
when "001100100100001" => rgb <= "000000";
when "001100100100010" => rgb <= "000000";
when "001100100100011" => rgb <= "000000";
when "001100100100100" => rgb <= "000000";
when "001100100100101" => rgb <= "000000";
when "001100100100110" => rgb <= "000000";
when "001100100101001" => rgb <= "000000";
when "001100100101010" => rgb <= "000000";
when "001100100101011" => rgb <= "000000";
when "001100100101100" => rgb <= "000000";
when "001100100101101" => rgb <= "000000";
when "001100100101110" => rgb <= "000000";
when "001100100101111" => rgb <= "000000";
when "001100100110010" => rgb <= "000000";
when "001100100110011" => rgb <= "000000";
when "001100100110100" => rgb <= "000000";
when "001100100110101" => rgb <= "000000";
when "001100100110110" => rgb <= "000000";
when "001100100110111" => rgb <= "000000";
when "001100100111000" => rgb <= "000000";
when "001100100111001" => rgb <= "000000";
when "001100100111010" => rgb <= "000000";
when "001100100111011" => rgb <= "000000";
when "001100100111100" => rgb <= "000000";
when "001100100111110" => rgb <= "000000";
when "001100100111111" => rgb <= "000000";
when "001100101000000" => rgb <= "000000";
when "001100101000001" => rgb <= "000000";
when "001100101000010" => rgb <= "000000";
when "001100101000011" => rgb <= "000000";
when "001100101000100" => rgb <= "000000";
when "001100101001000" => rgb <= "000000";
when "001100101001001" => rgb <= "000000";
when "001100101001010" => rgb <= "000000";
when "001100101001011" => rgb <= "000000";
when "001100101001100" => rgb <= "000000";
when "001100101001101" => rgb <= "000000";
when "001100101001110" => rgb <= "000000";
when "001100101011011" => rgb <= "000000";
when "001100101011100" => rgb <= "000000";
when "001100101011101" => rgb <= "000000";
when "001100101011110" => rgb <= "000000";
when "001100101011111" => rgb <= "000000";
when "001100101100000" => rgb <= "000000";
when "001100101100001" => rgb <= "000000";
when "001100101100010" => rgb <= "000000";
when "001100101100011" => rgb <= "000000";
when "001100101100100" => rgb <= "000000";
when "001100101100101" => rgb <= "000000";
when "001100101100110" => rgb <= "000000";
when "001100101100111" => rgb <= "000000";
when "001100101101000" => rgb <= "000000";
when "001100101101001" => rgb <= "000000";
when "001100101101010" => rgb <= "000000";
when "001100101101011" => rgb <= "000000";
when "001100101101100" => rgb <= "000000";
when "001100101101101" => rgb <= "000000";
when "001100101110000" => rgb <= "000000";
when "001100101110001" => rgb <= "000000";
when "001100101110010" => rgb <= "000000";
when "001100101110011" => rgb <= "000000";
when "001100101110100" => rgb <= "000000";
when "001100101110101" => rgb <= "000000";
when "001100101110110" => rgb <= "000000";
when "001100101110111" => rgb <= "000000";
when "001100101111000" => rgb <= "000000";
when "001100101111001" => rgb <= "000000";
when "001100101111010" => rgb <= "000000";
when "001100101111101" => rgb <= "000000";
when "001100101111110" => rgb <= "000000";
when "001100101111111" => rgb <= "000000";
when "001100110000000" => rgb <= "000000";
when "001100110000001" => rgb <= "000000";
when "001100110000010" => rgb <= "000000";
when "001100110000011" => rgb <= "000000";
when "001100110000100" => rgb <= "000000";
when "001100110000101" => rgb <= "000000";
when "001100110000110" => rgb <= "000000";
when "001100110000111" => rgb <= "000000";
when "001100110001000" => rgb <= "000000";
when "001100110001001" => rgb <= "000000";
when "001100110001010" => rgb <= "000000";
when "001100110001011" => rgb <= "000000";
when "001100110001100" => rgb <= "000000";
when "001100110001101" => rgb <= "000000";
when "001100110001110" => rgb <= "000000";
when "001100110001111" => rgb <= "000000";
when "001100110010000" => rgb <= "000000";
when "001100110010001" => rgb <= "000000";
when "001101000010001" => rgb <= "000000";
when "001101000010010" => rgb <= "000000";
when "001101000010011" => rgb <= "000000";
when "001101000010100" => rgb <= "000000";
when "001101000010101" => rgb <= "000000";
when "001101000010110" => rgb <= "000000";
when "001101000010111" => rgb <= "000000";
when "001101000011000" => rgb <= "000000";
when "001101000011001" => rgb <= "000000";
when "001101000011010" => rgb <= "000000";
when "001101000100001" => rgb <= "000000";
when "001101000100010" => rgb <= "000000";
when "001101000100011" => rgb <= "000000";
when "001101000100100" => rgb <= "000000";
when "001101000100101" => rgb <= "000000";
when "001101000100110" => rgb <= "000000";
when "001101000101010" => rgb <= "000000";
when "001101000101011" => rgb <= "000000";
when "001101000101100" => rgb <= "000000";
when "001101000101101" => rgb <= "000000";
when "001101000101110" => rgb <= "000000";
when "001101000101111" => rgb <= "000000";
when "001101000110011" => rgb <= "000000";
when "001101000110100" => rgb <= "000000";
when "001101000110101" => rgb <= "000000";
when "001101000110110" => rgb <= "000000";
when "001101000110111" => rgb <= "000000";
when "001101000111001" => rgb <= "000000";
when "001101000111010" => rgb <= "000000";
when "001101000111011" => rgb <= "000000";
when "001101000111100" => rgb <= "000000";
when "001101001000000" => rgb <= "000000";
when "001101001000001" => rgb <= "000000";
when "001101001000010" => rgb <= "000000";
when "001101001000011" => rgb <= "000000";
when "001101001000100" => rgb <= "000000";
when "001101001001001" => rgb <= "000000";
when "001101001001010" => rgb <= "000000";
when "001101001001011" => rgb <= "000000";
when "001101001001100" => rgb <= "000000";
when "001101001001101" => rgb <= "000000";
when "001101001001110" => rgb <= "000000";
when "001101001011011" => rgb <= "000000";
when "001101001011100" => rgb <= "000000";
when "001101001011101" => rgb <= "000000";
when "001101001011110" => rgb <= "000000";
when "001101001011111" => rgb <= "000000";
when "001101001100000" => rgb <= "000000";
when "001101001100001" => rgb <= "000000";
when "001101001100010" => rgb <= "000000";
when "001101001100011" => rgb <= "000000";
when "001101001100100" => rgb <= "000000";
when "001101001100101" => rgb <= "000000";
when "001101001100110" => rgb <= "000000";
when "001101001100111" => rgb <= "000000";
when "001101001101001" => rgb <= "000000";
when "001101001101010" => rgb <= "000000";
when "001101001101011" => rgb <= "000000";
when "001101001101100" => rgb <= "000000";
when "001101001101101" => rgb <= "000000";
when "001101001110001" => rgb <= "000000";
when "001101001110010" => rgb <= "000000";
when "001101001110011" => rgb <= "000000";
when "001101001110100" => rgb <= "000000";
when "001101001110101" => rgb <= "000000";
when "001101001110111" => rgb <= "000000";
when "001101001111000" => rgb <= "000000";
when "001101001111001" => rgb <= "000000";
when "001101001111010" => rgb <= "000000";
when "001101010000000" => rgb <= "000000";
when "001101010000001" => rgb <= "000000";
when "001101010000010" => rgb <= "000000";
when "001101010000011" => rgb <= "000000";
when "001101010000100" => rgb <= "000000";
when "001101010000110" => rgb <= "000000";
when "001101010000111" => rgb <= "000000";
when "001101010001000" => rgb <= "000000";
when "001101010001001" => rgb <= "000000";
when "001101010001010" => rgb <= "000000";
when "001101010001011" => rgb <= "000000";
when "001101010001100" => rgb <= "000000";
when "001101010001101" => rgb <= "000000";
when "001101010001110" => rgb <= "000000";
when "001101010001111" => rgb <= "000000";
when "001101010010000" => rgb <= "000000";
when "001101010010001" => rgb <= "000000";
when "001101100010001" => rgb <= "000000";
when "001101100010010" => rgb <= "000000";
when "001101100010011" => rgb <= "000000";
when "001101100010100" => rgb <= "000000";
when "001101100010101" => rgb <= "000000";
when "001101100010110" => rgb <= "000000";
when "001101100010111" => rgb <= "000000";
when "001101100011000" => rgb <= "000000";
when "001101100011001" => rgb <= "000000";
when "001101100011010" => rgb <= "000000";
when "001101100100001" => rgb <= "000000";
when "001101100100010" => rgb <= "000000";
when "001101100100011" => rgb <= "000000";
when "001101100100100" => rgb <= "000000";
when "001101100100101" => rgb <= "000000";
when "001101100100110" => rgb <= "000000";
when "001101100101010" => rgb <= "000000";
when "001101100101011" => rgb <= "000000";
when "001101100101100" => rgb <= "000000";
when "001101100101101" => rgb <= "000000";
when "001101100101110" => rgb <= "000000";
when "001101100101111" => rgb <= "000000";
when "001101100110011" => rgb <= "000000";
when "001101100110100" => rgb <= "000000";
when "001101100110101" => rgb <= "000000";
when "001101100110110" => rgb <= "000000";
when "001101100110111" => rgb <= "000000";
when "001101100111001" => rgb <= "000000";
when "001101100111010" => rgb <= "000000";
when "001101100111011" => rgb <= "000000";
when "001101100111100" => rgb <= "000000";
when "001101101000000" => rgb <= "000000";
when "001101101000001" => rgb <= "000000";
when "001101101000010" => rgb <= "000000";
when "001101101000011" => rgb <= "000000";
when "001101101000100" => rgb <= "000000";
when "001101101001001" => rgb <= "000000";
when "001101101001010" => rgb <= "000000";
when "001101101001011" => rgb <= "000000";
when "001101101001100" => rgb <= "000000";
when "001101101001101" => rgb <= "000000";
when "001101101001110" => rgb <= "000000";
when "001101101011100" => rgb <= "000000";
when "001101101011101" => rgb <= "000000";
when "001101101011110" => rgb <= "000000";
when "001101101011111" => rgb <= "000000";
when "001101101100000" => rgb <= "000000";
when "001101101100001" => rgb <= "000000";
when "001101101100010" => rgb <= "000000";
when "001101101100011" => rgb <= "000000";
when "001101101100100" => rgb <= "000000";
when "001101101100101" => rgb <= "000000";
when "001101101100110" => rgb <= "000000";
when "001101101100111" => rgb <= "000000";
when "001101101101001" => rgb <= "000000";
when "001101101101010" => rgb <= "000000";
when "001101101101011" => rgb <= "000000";
when "001101101101100" => rgb <= "000000";
when "001101101101101" => rgb <= "000000";
when "001101101110001" => rgb <= "000000";
when "001101101110010" => rgb <= "000000";
when "001101101110011" => rgb <= "000000";
when "001101101110100" => rgb <= "000000";
when "001101101110101" => rgb <= "000000";
when "001101101110111" => rgb <= "000000";
when "001101101111000" => rgb <= "000000";
when "001101101111001" => rgb <= "000000";
when "001101101111010" => rgb <= "000000";
when "001101110000000" => rgb <= "000000";
when "001101110000001" => rgb <= "000000";
when "001101110000010" => rgb <= "000000";
when "001101110000011" => rgb <= "000000";
when "001101110000100" => rgb <= "000000";
when "001101110000110" => rgb <= "000000";
when "001101110000111" => rgb <= "000000";
when "001101110001000" => rgb <= "000000";
when "001101110001001" => rgb <= "000000";
when "001101110001010" => rgb <= "000000";
when "001101110001011" => rgb <= "000000";
when "001101110001100" => rgb <= "000000";
when "001101110001101" => rgb <= "000000";
when "001101110001110" => rgb <= "000000";
when "001101110001111" => rgb <= "000000";
when "001101110010000" => rgb <= "000000";
when "001101110010001" => rgb <= "000000";
when "010100101001001" => rgb <= "000000";
when "010100101001010" => rgb <= "000000";
when "010100101001011" => rgb <= "000000";
when "010100101001101" => rgb <= "000000";
when "010100101010001" => rgb <= "000000";
when "010100101010010" => rgb <= "000000";
when "010100101010011" => rgb <= "000000";
when "010100101010101" => rgb <= "000000";
when "010100101010111" => rgb <= "000000";
when "010101001001001" => rgb <= "000000";
when "010101001001011" => rgb <= "000000";
when "010101001001101" => rgb <= "000000";
when "010101001010001" => rgb <= "000000";
when "010101001010011" => rgb <= "000000";
when "010101001010101" => rgb <= "000000";
when "010101001010111" => rgb <= "000000";
when "010101101001001" => rgb <= "000000";
when "010101101001010" => rgb <= "000000";
when "010101101001011" => rgb <= "000000";
when "010101101001101" => rgb <= "000000";
when "010101101010001" => rgb <= "000000";
when "010101101010010" => rgb <= "000000";
when "010101101010011" => rgb <= "000000";
when "010101101010101" => rgb <= "000000";
when "010101101010111" => rgb <= "000000";
when "010110001001001" => rgb <= "000000";
when "010110001001101" => rgb <= "000000";
when "010110001010001" => rgb <= "000000";
when "010110001010011" => rgb <= "000000";
when "010110001010110" => rgb <= "000000";
when "010110101001001" => rgb <= "000000";
when "010110101001101" => rgb <= "000000";
when "010110101001110" => rgb <= "000000";
when "010110101001111" => rgb <= "000000";
when "010110101010001" => rgb <= "000000";
when "010110101010011" => rgb <= "000000";
when "010110101010110" => rgb <= "000000";
                when others => rgb <= "111111"; --will update l8r
            end case;
        end if;
    end process; 
	addressOut <= address;
end;  