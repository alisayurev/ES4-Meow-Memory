library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;


entity two is 
port(
    clk : in std_logic;
	address : in unsigned (14 downto 0); 
    rgb : out unsigned(5 downto 0)
);
end two;


architecture synth of two is 

signal addressOut : unsigned(14 downto 0); 

begin
    process (clk) is begin
        if rising_edge(clk) then
            case addressOut is
			when "000011000111000" => rgb <= "000000";

when "000011000111001" => rgb <= "000000";

when "000011000111010" => rgb <= "000000";

when "000011000111011" => rgb <= "000000";

when "000011000111100" => rgb <= "000000";

when "000011000111101" => rgb <= "000000";

when "000011000111110" => rgb <= "000000";

when "000011000111111" => rgb <= "000000";

when "000011001000000" => rgb <= "000000";

when "000011001000001" => rgb <= "000000";

when "000011001000010" => rgb <= "000000";

when "000011001000011" => rgb <= "000000";

when "000011001000100" => rgb <= "000000";

when "000011001000101" => rgb <= "000000";

when "000011001000110" => rgb <= "000000";

when "000011001000111" => rgb <= "000000";

when "000011001001000" => rgb <= "000000";

when "000011001001001" => rgb <= "000000";

when "000011001001010" => rgb <= "000000";

when "000011001001011" => rgb <= "000000";

when "000011001001100" => rgb <= "000000";

when "000011001001101" => rgb <= "000000";

when "000011001001110" => rgb <= "000000";

when "000011001001111" => rgb <= "000000";

when "000011001010000" => rgb <= "000000";

when "000011001010001" => rgb <= "000000";

when "000011001010010" => rgb <= "000000";

when "000011001010011" => rgb <= "000000";

when "000011001010100" => rgb <= "000000";

when "000011001010101" => rgb <= "000000";

when "000011001010110" => rgb <= "000000";

when "000011001010111" => rgb <= "000000";

when "000011001011000" => rgb <= "000000";

when "000011001011001" => rgb <= "000000";

when "000011001011010" => rgb <= "000000";

when "000011001011011" => rgb <= "000000";

when "000011001011100" => rgb <= "000000";

when "000011001011101" => rgb <= "000000";

when "000011001011110" => rgb <= "000000";

when "000011001011111" => rgb <= "000000";

when "000011001100000" => rgb <= "000000";

when "000011001100001" => rgb <= "000000";

when "000011001100010" => rgb <= "000000";

when "000011001100011" => rgb <= "000000";

when "000011001100100" => rgb <= "000000";

when "000011001100101" => rgb <= "000000";

when "000011001100110" => rgb <= "000000";

when "000011001100111" => rgb <= "000000";

when "000011100111000" => rgb <= "000000";

when "000011100111001" => rgb <= "100110";

when "000011100111010" => rgb <= "100110";

when "000011100111011" => rgb <= "100110";

when "000011100111100" => rgb <= "100110";

when "000011100111101" => rgb <= "100110";

when "000011100111110" => rgb <= "100110";

when "000011100111111" => rgb <= "100110";

when "000011101000000" => rgb <= "100110";

when "000011101000001" => rgb <= "100110";

when "000011101000010" => rgb <= "100110";

when "000011101000011" => rgb <= "100110";

when "000011101000100" => rgb <= "100110";

when "000011101000101" => rgb <= "100110";

when "000011101000110" => rgb <= "100110";

when "000011101000111" => rgb <= "100110";

when "000011101001000" => rgb <= "100110";

when "000011101001001" => rgb <= "100110";

when "000011101001010" => rgb <= "100110";

when "000011101001011" => rgb <= "100110";

when "000011101001100" => rgb <= "100110";

when "000011101001101" => rgb <= "100110";

when "000011101001110" => rgb <= "100110";

when "000011101001111" => rgb <= "100110";

when "000011101010000" => rgb <= "100110";

when "000011101010001" => rgb <= "100110";

when "000011101010010" => rgb <= "100110";

when "000011101010011" => rgb <= "100110";

when "000011101010100" => rgb <= "100110";

when "000011101010101" => rgb <= "100110";

when "000011101010110" => rgb <= "100110";

when "000011101010111" => rgb <= "100110";

when "000011101011000" => rgb <= "100110";

when "000011101011001" => rgb <= "100110";

when "000011101011010" => rgb <= "100110";

when "000011101011011" => rgb <= "100110";

when "000011101011100" => rgb <= "100110";

when "000011101011101" => rgb <= "100110";

when "000011101011110" => rgb <= "100110";

when "000011101011111" => rgb <= "100110";

when "000011101100000" => rgb <= "100110";

when "000011101100001" => rgb <= "100110";

when "000011101100010" => rgb <= "100110";

when "000011101100011" => rgb <= "100110";

when "000011101100100" => rgb <= "100110";

when "000011101100101" => rgb <= "100110";

when "000011101100110" => rgb <= "100110";

when "000011101100111" => rgb <= "000000";

when "000100000111000" => rgb <= "000000";

when "000100000111001" => rgb <= "100110";

when "000100000111010" => rgb <= "100110";

when "000100000111011" => rgb <= "100110";

when "000100000111100" => rgb <= "100110";

when "000100000111101" => rgb <= "100110";

when "000100000111110" => rgb <= "100110";

when "000100000111111" => rgb <= "100110";

when "000100001000000" => rgb <= "100110";

when "000100001000001" => rgb <= "100110";

when "000100001000010" => rgb <= "100110";

when "000100001000011" => rgb <= "100110";

when "000100001000100" => rgb <= "100110";

when "000100001000101" => rgb <= "100110";

when "000100001000110" => rgb <= "100110";

when "000100001000111" => rgb <= "100110";

when "000100001001000" => rgb <= "100110";

when "000100001001001" => rgb <= "100110";

when "000100001001010" => rgb <= "100110";

when "000100001001011" => rgb <= "100110";

when "000100001001100" => rgb <= "100110";

when "000100001001101" => rgb <= "100110";

when "000100001001110" => rgb <= "100110";

when "000100001001111" => rgb <= "100110";

when "000100001010000" => rgb <= "100110";

when "000100001010001" => rgb <= "100110";

when "000100001010010" => rgb <= "100110";

when "000100001010011" => rgb <= "100110";

when "000100001010100" => rgb <= "100110";

when "000100001010101" => rgb <= "100110";

when "000100001010110" => rgb <= "100110";

when "000100001010111" => rgb <= "100110";

when "000100001011000" => rgb <= "100110";

when "000100001011001" => rgb <= "100110";

when "000100001011010" => rgb <= "100110";

when "000100001011011" => rgb <= "100110";

when "000100001011100" => rgb <= "100110";

when "000100001011101" => rgb <= "100110";

when "000100001011110" => rgb <= "100110";

when "000100001011111" => rgb <= "100110";

when "000100001100000" => rgb <= "100110";

when "000100001100001" => rgb <= "100110";

when "000100001100010" => rgb <= "100110";

when "000100001100011" => rgb <= "100110";

when "000100001100100" => rgb <= "100110";

when "000100001100101" => rgb <= "100110";

when "000100001100110" => rgb <= "100110";

when "000100001100111" => rgb <= "000000";

when "000100100111000" => rgb <= "000000";

when "000100100111001" => rgb <= "100110";

when "000100100111010" => rgb <= "100110";

when "000100100111011" => rgb <= "100110";

when "000100100111100" => rgb <= "100110";

when "000100100111101" => rgb <= "100110";

when "000100100111110" => rgb <= "100110";

when "000100100111111" => rgb <= "100110";

when "000100101000000" => rgb <= "100110";

when "000100101000001" => rgb <= "100110";

when "000100101000010" => rgb <= "100110";

when "000100101000011" => rgb <= "100110";

when "000100101000100" => rgb <= "100110";

when "000100101000101" => rgb <= "100110";

when "000100101000110" => rgb <= "100110";

when "000100101000111" => rgb <= "100110";

when "000100101001000" => rgb <= "100110";

when "000100101001001" => rgb <= "100110";

when "000100101001010" => rgb <= "100110";

when "000100101001011" => rgb <= "100110";

when "000100101001100" => rgb <= "100110";

when "000100101001101" => rgb <= "100110";

when "000100101001110" => rgb <= "100110";

when "000100101001111" => rgb <= "100110";

when "000100101010000" => rgb <= "100110";

when "000100101010001" => rgb <= "100110";

when "000100101010010" => rgb <= "100110";

when "000100101010011" => rgb <= "100110";

when "000100101010100" => rgb <= "100110";

when "000100101010101" => rgb <= "100110";

when "000100101010110" => rgb <= "100110";

when "000100101010111" => rgb <= "100110";

when "000100101011000" => rgb <= "100110";

when "000100101011001" => rgb <= "100110";

when "000100101011010" => rgb <= "100110";

when "000100101011011" => rgb <= "100110";

when "000100101011100" => rgb <= "100110";

when "000100101011101" => rgb <= "100110";

when "000100101011110" => rgb <= "100110";

when "000100101011111" => rgb <= "100110";

when "000100101100000" => rgb <= "100110";

when "000100101100001" => rgb <= "100110";

when "000100101100010" => rgb <= "100110";

when "000100101100011" => rgb <= "100110";

when "000100101100100" => rgb <= "100110";

when "000100101100101" => rgb <= "100110";

when "000100101100110" => rgb <= "100110";

when "000100101100111" => rgb <= "000000";

when "000101000111000" => rgb <= "000000";

when "000101000111001" => rgb <= "100110";

when "000101000111010" => rgb <= "100110";

when "000101000111011" => rgb <= "100110";

when "000101000111100" => rgb <= "100110";

when "000101000111101" => rgb <= "100110";

when "000101000111110" => rgb <= "100110";

when "000101000111111" => rgb <= "100110";

when "000101001000000" => rgb <= "100110";

when "000101001000001" => rgb <= "100110";

when "000101001000010" => rgb <= "100110";

when "000101001000011" => rgb <= "100110";

when "000101001000100" => rgb <= "100110";

when "000101001000101" => rgb <= "100110";

when "000101001000110" => rgb <= "100110";

when "000101001000111" => rgb <= "100110";

when "000101001001000" => rgb <= "100110";

when "000101001001001" => rgb <= "100110";

when "000101001001010" => rgb <= "100110";

when "000101001001011" => rgb <= "100110";

when "000101001001100" => rgb <= "100110";

when "000101001001101" => rgb <= "100110";

when "000101001001110" => rgb <= "100110";

when "000101001001111" => rgb <= "100110";

when "000101001010000" => rgb <= "100110";

when "000101001010001" => rgb <= "100110";

when "000101001010010" => rgb <= "100110";

when "000101001010011" => rgb <= "100110";

when "000101001010100" => rgb <= "100110";

when "000101001010101" => rgb <= "100110";

when "000101001010110" => rgb <= "100110";

when "000101001010111" => rgb <= "100110";

when "000101001011000" => rgb <= "100110";

when "000101001011001" => rgb <= "100110";

when "000101001011010" => rgb <= "100110";

when "000101001011011" => rgb <= "100110";

when "000101001011100" => rgb <= "100110";

when "000101001011101" => rgb <= "100110";

when "000101001011110" => rgb <= "100110";

when "000101001011111" => rgb <= "100110";

when "000101001100000" => rgb <= "100110";

when "000101001100001" => rgb <= "100110";

when "000101001100010" => rgb <= "100110";

when "000101001100011" => rgb <= "100110";

when "000101001100100" => rgb <= "100110";

when "000101001100101" => rgb <= "100110";

when "000101001100110" => rgb <= "100110";

when "000101001100111" => rgb <= "000000";

when "000101100111000" => rgb <= "000000";

when "000101100111001" => rgb <= "100110";

when "000101100111010" => rgb <= "100110";

when "000101100111011" => rgb <= "100110";

when "000101100111100" => rgb <= "100110";

when "000101100111101" => rgb <= "100110";

when "000101100111110" => rgb <= "100110";

when "000101100111111" => rgb <= "100110";

when "000101101000000" => rgb <= "100110";

when "000101101000001" => rgb <= "100110";

when "000101101000010" => rgb <= "100110";

when "000101101000011" => rgb <= "100110";

when "000101101000100" => rgb <= "100110";

when "000101101000101" => rgb <= "100110";

when "000101101000110" => rgb <= "100110";

when "000101101000111" => rgb <= "100110";

when "000101101001000" => rgb <= "100110";

when "000101101001001" => rgb <= "100110";

when "000101101001010" => rgb <= "100110";

when "000101101001011" => rgb <= "100110";

when "000101101001100" => rgb <= "100110";

when "000101101001101" => rgb <= "100110";

when "000101101001110" => rgb <= "100110";

when "000101101001111" => rgb <= "100110";

when "000101101010000" => rgb <= "100110";

when "000101101010001" => rgb <= "100110";

when "000101101010010" => rgb <= "100110";

when "000101101010011" => rgb <= "100110";

when "000101101010100" => rgb <= "100110";

when "000101101010101" => rgb <= "100110";

when "000101101010110" => rgb <= "100110";

when "000101101010111" => rgb <= "100110";

when "000101101011000" => rgb <= "100110";

when "000101101011001" => rgb <= "100110";

when "000101101011010" => rgb <= "100110";

when "000101101011011" => rgb <= "100110";

when "000101101011100" => rgb <= "100110";

when "000101101011101" => rgb <= "100110";

when "000101101011110" => rgb <= "100110";

when "000101101011111" => rgb <= "100110";

when "000101101100000" => rgb <= "100110";

when "000101101100001" => rgb <= "100110";

when "000101101100010" => rgb <= "100110";

when "000101101100011" => rgb <= "100110";

when "000101101100100" => rgb <= "100110";

when "000101101100101" => rgb <= "100110";

when "000101101100110" => rgb <= "100110";

when "000101101100111" => rgb <= "000000";

when "000110000111000" => rgb <= "000000";

when "000110000111001" => rgb <= "100110";

when "000110000111010" => rgb <= "100110";

when "000110000111011" => rgb <= "100110";

when "000110000111100" => rgb <= "100110";

when "000110000111101" => rgb <= "100110";

when "000110000111110" => rgb <= "100110";

when "000110000111111" => rgb <= "100110";

when "000110001000000" => rgb <= "100110";

when "000110001000001" => rgb <= "100110";

when "000110001000010" => rgb <= "100110";

when "000110001000011" => rgb <= "100110";

when "000110001000100" => rgb <= "100110";

when "000110001000101" => rgb <= "100110";

when "000110001000110" => rgb <= "100110";

when "000110001000111" => rgb <= "100110";

when "000110001001000" => rgb <= "100110";

when "000110001001001" => rgb <= "100110";

when "000110001001010" => rgb <= "100110";

when "000110001001011" => rgb <= "100110";

when "000110001001100" => rgb <= "100110";

when "000110001001101" => rgb <= "100110";

when "000110001001110" => rgb <= "100110";

when "000110001001111" => rgb <= "100110";

when "000110001010000" => rgb <= "100110";

when "000110001010001" => rgb <= "100110";

when "000110001010010" => rgb <= "100110";

when "000110001010011" => rgb <= "100110";

when "000110001010100" => rgb <= "100110";

when "000110001010101" => rgb <= "100110";

when "000110001010110" => rgb <= "100110";

when "000110001010111" => rgb <= "100110";

when "000110001011000" => rgb <= "100110";

when "000110001011001" => rgb <= "100110";

when "000110001011010" => rgb <= "100110";

when "000110001011011" => rgb <= "100110";

when "000110001011100" => rgb <= "100110";

when "000110001011101" => rgb <= "100110";

when "000110001011110" => rgb <= "100110";

when "000110001011111" => rgb <= "100110";

when "000110001100000" => rgb <= "100110";

when "000110001100001" => rgb <= "100110";

when "000110001100010" => rgb <= "100110";

when "000110001100011" => rgb <= "100110";

when "000110001100100" => rgb <= "100110";

when "000110001100101" => rgb <= "100110";

when "000110001100110" => rgb <= "100110";

when "000110001100111" => rgb <= "000000";

when "000110100111000" => rgb <= "000000";

when "000110100111001" => rgb <= "100110";

when "000110100111010" => rgb <= "100110";

when "000110100111011" => rgb <= "100110";

when "000110100111100" => rgb <= "100110";

when "000110100111101" => rgb <= "100110";

when "000110100111110" => rgb <= "100110";

when "000110100111111" => rgb <= "000000";

when "000110101000000" => rgb <= "000000";

when "000110101000001" => rgb <= "000000";

when "000110101000010" => rgb <= "000000";

when "000110101000011" => rgb <= "000000";

when "000110101000100" => rgb <= "000000";

when "000110101000101" => rgb <= "000000";

when "000110101000110" => rgb <= "000000";

when "000110101000111" => rgb <= "000000";

when "000110101001000" => rgb <= "000000";

when "000110101001001" => rgb <= "000000";

when "000110101001010" => rgb <= "000000";

when "000110101001011" => rgb <= "000000";

when "000110101001100" => rgb <= "000000";

when "000110101001101" => rgb <= "000000";

when "000110101001110" => rgb <= "000000";

when "000110101001111" => rgb <= "000000";

when "000110101010000" => rgb <= "000000";

when "000110101010001" => rgb <= "000000";

when "000110101010010" => rgb <= "000000";

when "000110101010011" => rgb <= "000000";

when "000110101010100" => rgb <= "000000";

when "000110101010101" => rgb <= "000000";

when "000110101010110" => rgb <= "000000";

when "000110101010111" => rgb <= "000000";

when "000110101011000" => rgb <= "000000";

when "000110101011001" => rgb <= "000000";

when "000110101011010" => rgb <= "000000";

when "000110101011011" => rgb <= "000000";

when "000110101011100" => rgb <= "000000";

when "000110101011101" => rgb <= "000000";

when "000110101011110" => rgb <= "000000";

when "000110101011111" => rgb <= "100110";

when "000110101100000" => rgb <= "100110";

when "000110101100001" => rgb <= "100110";

when "000110101100010" => rgb <= "100110";

when "000110101100011" => rgb <= "100110";

when "000110101100100" => rgb <= "100110";

when "000110101100101" => rgb <= "100110";

when "000110101100110" => rgb <= "100110";

when "000110101100111" => rgb <= "000000";

when "000111000111000" => rgb <= "000000";

when "000111000111001" => rgb <= "100110";

when "000111000111010" => rgb <= "100110";

when "000111000111011" => rgb <= "100110";

when "000111000111100" => rgb <= "100110";

when "000111000111101" => rgb <= "100110";

when "000111000111110" => rgb <= "100110";

when "000111000111111" => rgb <= "000000";

when "000111001011110" => rgb <= "000000";

when "000111001011111" => rgb <= "100110";

when "000111001100000" => rgb <= "100110";

when "000111001100001" => rgb <= "100110";

when "000111001100010" => rgb <= "100110";

when "000111001100011" => rgb <= "100110";

when "000111001100100" => rgb <= "100110";

when "000111001100101" => rgb <= "100110";

when "000111001100110" => rgb <= "100110";

when "000111001100111" => rgb <= "000000";

when "000111100111000" => rgb <= "000000";

when "000111100111001" => rgb <= "100110";

when "000111100111010" => rgb <= "100110";

when "000111100111011" => rgb <= "100110";

when "000111100111100" => rgb <= "100110";

when "000111100111101" => rgb <= "100110";

when "000111100111110" => rgb <= "100110";

when "000111100111111" => rgb <= "000000";

when "000111101011110" => rgb <= "000000";

when "000111101011111" => rgb <= "100110";

when "000111101100000" => rgb <= "100110";

when "000111101100001" => rgb <= "100110";

when "000111101100010" => rgb <= "100110";

when "000111101100011" => rgb <= "100110";

when "000111101100100" => rgb <= "100110";

when "000111101100101" => rgb <= "100110";

when "000111101100110" => rgb <= "100110";

when "000111101100111" => rgb <= "000000";

when "001000000111000" => rgb <= "000000";

when "001000000111001" => rgb <= "100110";

when "001000000111010" => rgb <= "100110";

when "001000000111011" => rgb <= "100110";

when "001000000111100" => rgb <= "100110";

when "001000000111101" => rgb <= "100110";

when "001000000111110" => rgb <= "100110";

when "001000000111111" => rgb <= "000000";

when "001000001011110" => rgb <= "000000";

when "001000001011111" => rgb <= "100110";

when "001000001100000" => rgb <= "100110";

when "001000001100001" => rgb <= "100110";

when "001000001100010" => rgb <= "100110";

when "001000001100011" => rgb <= "100110";

when "001000001100100" => rgb <= "100110";

when "001000001100101" => rgb <= "100110";

when "001000001100110" => rgb <= "100110";

when "001000001100111" => rgb <= "000000";

when "001000100111000" => rgb <= "000000";

when "001000100111001" => rgb <= "100110";

when "001000100111010" => rgb <= "100110";

when "001000100111011" => rgb <= "100110";

when "001000100111100" => rgb <= "100110";

when "001000100111101" => rgb <= "100110";

when "001000100111110" => rgb <= "100110";

when "001000100111111" => rgb <= "000000";

when "001000101011110" => rgb <= "000000";

when "001000101011111" => rgb <= "100110";

when "001000101100000" => rgb <= "100110";

when "001000101100001" => rgb <= "100110";

when "001000101100010" => rgb <= "100110";

when "001000101100011" => rgb <= "100110";

when "001000101100100" => rgb <= "100110";

when "001000101100101" => rgb <= "100110";

when "001000101100110" => rgb <= "100110";

when "001000101100111" => rgb <= "000000";

when "001001000111000" => rgb <= "000000";

when "001001000111001" => rgb <= "000000";

when "001001000111010" => rgb <= "000000";

when "001001000111011" => rgb <= "000000";

when "001001000111100" => rgb <= "000000";

when "001001000111101" => rgb <= "000000";

when "001001000111110" => rgb <= "000000";

when "001001000111111" => rgb <= "000000";

when "001001001011110" => rgb <= "000000";

when "001001001011111" => rgb <= "100110";

when "001001001100000" => rgb <= "100110";

when "001001001100001" => rgb <= "100110";

when "001001001100010" => rgb <= "100110";

when "001001001100011" => rgb <= "100110";

when "001001001100100" => rgb <= "100110";

when "001001001100101" => rgb <= "100110";

when "001001001100110" => rgb <= "100110";

when "001001001100111" => rgb <= "000000";

when "001001101011110" => rgb <= "000000";

when "001001101011111" => rgb <= "100110";

when "001001101100000" => rgb <= "100110";

when "001001101100001" => rgb <= "100110";

when "001001101100010" => rgb <= "100110";

when "001001101100011" => rgb <= "100110";

when "001001101100100" => rgb <= "100110";

when "001001101100101" => rgb <= "100110";

when "001001101100110" => rgb <= "100110";

when "001001101100111" => rgb <= "000000";

when "001010001011110" => rgb <= "000000";

when "001010001011111" => rgb <= "100110";

when "001010001100000" => rgb <= "100110";

when "001010001100001" => rgb <= "100110";

when "001010001100010" => rgb <= "100110";

when "001010001100011" => rgb <= "100110";

when "001010001100100" => rgb <= "100110";

when "001010001100101" => rgb <= "100110";

when "001010001100110" => rgb <= "100110";

when "001010001100111" => rgb <= "000000";

when "001010101011110" => rgb <= "000000";

when "001010101011111" => rgb <= "100110";

when "001010101100000" => rgb <= "100110";

when "001010101100001" => rgb <= "100110";

when "001010101100010" => rgb <= "100110";

when "001010101100011" => rgb <= "100110";

when "001010101100100" => rgb <= "100110";

when "001010101100101" => rgb <= "100110";

when "001010101100110" => rgb <= "100110";

when "001010101100111" => rgb <= "000000";

when "001011001011110" => rgb <= "000000";

when "001011001011111" => rgb <= "100110";

when "001011001100000" => rgb <= "100110";

when "001011001100001" => rgb <= "100110";

when "001011001100010" => rgb <= "100110";

when "001011001100011" => rgb <= "100110";

when "001011001100100" => rgb <= "100110";

when "001011001100101" => rgb <= "100110";

when "001011001100110" => rgb <= "100110";

when "001011001100111" => rgb <= "000000";

when "001011101011110" => rgb <= "000000";

when "001011101011111" => rgb <= "100110";

when "001011101100000" => rgb <= "100110";

when "001011101100001" => rgb <= "100110";

when "001011101100010" => rgb <= "100110";

when "001011101100011" => rgb <= "100110";

when "001011101100100" => rgb <= "100110";

when "001011101100101" => rgb <= "100110";

when "001011101100110" => rgb <= "100110";

when "001011101100111" => rgb <= "000000";

when "001100001011110" => rgb <= "000000";

when "001100001011111" => rgb <= "100110";

when "001100001100000" => rgb <= "100110";

when "001100001100001" => rgb <= "100110";

when "001100001100010" => rgb <= "100110";

when "001100001100011" => rgb <= "100110";

when "001100001100100" => rgb <= "100110";

when "001100001100101" => rgb <= "100110";

when "001100001100110" => rgb <= "100110";

when "001100001100111" => rgb <= "000000";

when "001100101011110" => rgb <= "000000";

when "001100101011111" => rgb <= "100110";

when "001100101100000" => rgb <= "100110";

when "001100101100001" => rgb <= "100110";

when "001100101100010" => rgb <= "100110";

when "001100101100011" => rgb <= "100110";

when "001100101100100" => rgb <= "100110";

when "001100101100101" => rgb <= "100110";

when "001100101100110" => rgb <= "100110";

when "001100101100111" => rgb <= "000000";

when "001101001011110" => rgb <= "000000";

when "001101001011111" => rgb <= "100110";

when "001101001100000" => rgb <= "100110";

when "001101001100001" => rgb <= "100110";

when "001101001100010" => rgb <= "100110";

when "001101001100011" => rgb <= "100110";

when "001101001100100" => rgb <= "100110";

when "001101001100101" => rgb <= "100110";

when "001101001100110" => rgb <= "100110";

when "001101001100111" => rgb <= "000000";

when "001101101011110" => rgb <= "000000";

when "001101101011111" => rgb <= "100110";

when "001101101100000" => rgb <= "100110";

when "001101101100001" => rgb <= "100110";

when "001101101100010" => rgb <= "100110";

when "001101101100011" => rgb <= "100110";

when "001101101100100" => rgb <= "100110";

when "001101101100101" => rgb <= "100110";

when "001101101100110" => rgb <= "100110";

when "001101101100111" => rgb <= "000000";

when "001110001011110" => rgb <= "000000";

when "001110001011111" => rgb <= "100110";

when "001110001100000" => rgb <= "100110";

when "001110001100001" => rgb <= "100110";

when "001110001100010" => rgb <= "100110";

when "001110001100011" => rgb <= "100110";

when "001110001100100" => rgb <= "100110";

when "001110001100101" => rgb <= "100110";

when "001110001100110" => rgb <= "100110";

when "001110001100111" => rgb <= "000000";

when "001110101011110" => rgb <= "000000";

when "001110101011111" => rgb <= "100110";

when "001110101100000" => rgb <= "100110";

when "001110101100001" => rgb <= "100110";

when "001110101100010" => rgb <= "100110";

when "001110101100011" => rgb <= "100110";

when "001110101100100" => rgb <= "100110";

when "001110101100101" => rgb <= "100110";

when "001110101100110" => rgb <= "100110";

when "001110101100111" => rgb <= "000000";

when "001111001011110" => rgb <= "000000";

when "001111001011111" => rgb <= "100110";

when "001111001100000" => rgb <= "100110";

when "001111001100001" => rgb <= "100110";

when "001111001100010" => rgb <= "100110";

when "001111001100011" => rgb <= "100110";

when "001111001100100" => rgb <= "100110";

when "001111001100101" => rgb <= "100110";

when "001111001100110" => rgb <= "100110";

when "001111001100111" => rgb <= "000000";

when "001111100111000" => rgb <= "000000";

when "001111100111001" => rgb <= "000000";

when "001111100111010" => rgb <= "000000";

when "001111100111011" => rgb <= "000000";

when "001111100111100" => rgb <= "000000";

when "001111100111101" => rgb <= "000000";

when "001111100111110" => rgb <= "000000";

when "001111100111111" => rgb <= "000000";

when "001111101000000" => rgb <= "000000";

when "001111101000001" => rgb <= "000000";

when "001111101000010" => rgb <= "000000";

when "001111101000011" => rgb <= "000000";

when "001111101000100" => rgb <= "000000";

when "001111101000101" => rgb <= "000000";

when "001111101000110" => rgb <= "000000";

when "001111101000111" => rgb <= "000000";

when "001111101001000" => rgb <= "000000";

when "001111101001001" => rgb <= "000000";

when "001111101001010" => rgb <= "000000";

when "001111101001011" => rgb <= "000000";

when "001111101001100" => rgb <= "000000";

when "001111101001101" => rgb <= "000000";

when "001111101001110" => rgb <= "000000";

when "001111101001111" => rgb <= "000000";

when "001111101010000" => rgb <= "000000";

when "001111101010001" => rgb <= "000000";

when "001111101010010" => rgb <= "000000";

when "001111101010011" => rgb <= "000000";

when "001111101010100" => rgb <= "000000";

when "001111101010101" => rgb <= "000000";

when "001111101010110" => rgb <= "000000";

when "001111101010111" => rgb <= "000000";

when "001111101011000" => rgb <= "000000";

when "001111101011001" => rgb <= "000000";

when "001111101011010" => rgb <= "000000";

when "001111101011011" => rgb <= "000000";

when "001111101011100" => rgb <= "000000";

when "001111101011101" => rgb <= "000000";

when "001111101011110" => rgb <= "000000";

when "001111101011111" => rgb <= "100110";

when "001111101100000" => rgb <= "100110";

when "001111101100001" => rgb <= "100110";

when "001111101100010" => rgb <= "100110";

when "001111101100011" => rgb <= "100110";

when "001111101100100" => rgb <= "100110";

when "001111101100101" => rgb <= "100110";

when "001111101100110" => rgb <= "100110";

when "001111101100111" => rgb <= "000000";

when "010000000111000" => rgb <= "000000";

when "010000000111001" => rgb <= "100110";

when "010000000111010" => rgb <= "100110";

when "010000000111011" => rgb <= "100110";

when "010000000111100" => rgb <= "100110";

when "010000000111101" => rgb <= "100110";

when "010000000111110" => rgb <= "100110";

when "010000000111111" => rgb <= "100110";

when "010000001000000" => rgb <= "100110";

when "010000001000001" => rgb <= "100110";

when "010000001000010" => rgb <= "100110";

when "010000001000011" => rgb <= "100110";

when "010000001000100" => rgb <= "100110";

when "010000001000101" => rgb <= "100110";

when "010000001000110" => rgb <= "100110";

when "010000001000111" => rgb <= "100110";

when "010000001001000" => rgb <= "100110";

when "010000001001001" => rgb <= "100110";

when "010000001001010" => rgb <= "100110";

when "010000001001011" => rgb <= "100110";

when "010000001001100" => rgb <= "100110";

when "010000001001101" => rgb <= "100110";

when "010000001001110" => rgb <= "100110";

when "010000001001111" => rgb <= "100110";

when "010000001010000" => rgb <= "100110";

when "010000001010001" => rgb <= "100110";

when "010000001010010" => rgb <= "100110";

when "010000001010011" => rgb <= "100110";

when "010000001010100" => rgb <= "100110";

when "010000001010101" => rgb <= "100110";

when "010000001010110" => rgb <= "100110";

when "010000001010111" => rgb <= "100110";

when "010000001011000" => rgb <= "100110";

when "010000001011001" => rgb <= "100110";

when "010000001011010" => rgb <= "100110";

when "010000001011011" => rgb <= "100110";

when "010000001011100" => rgb <= "100110";

when "010000001011101" => rgb <= "100110";

when "010000001011110" => rgb <= "100110";

when "010000001011111" => rgb <= "100110";

when "010000001100000" => rgb <= "100110";

when "010000001100001" => rgb <= "100110";

when "010000001100010" => rgb <= "100110";

when "010000001100011" => rgb <= "100110";

when "010000001100100" => rgb <= "100110";

when "010000001100101" => rgb <= "100110";

when "010000001100110" => rgb <= "100110";

when "010000001100111" => rgb <= "000000";

when "010000100111000" => rgb <= "000000";

when "010000100111001" => rgb <= "100110";

when "010000100111010" => rgb <= "100110";

when "010000100111011" => rgb <= "100110";

when "010000100111100" => rgb <= "100110";

when "010000100111101" => rgb <= "100110";

when "010000100111110" => rgb <= "100110";

when "010000100111111" => rgb <= "100110";

when "010000101000000" => rgb <= "100110";

when "010000101000001" => rgb <= "100110";

when "010000101000010" => rgb <= "100110";

when "010000101000011" => rgb <= "100110";

when "010000101000100" => rgb <= "100110";

when "010000101000101" => rgb <= "100110";

when "010000101000110" => rgb <= "100110";

when "010000101000111" => rgb <= "100110";

when "010000101001000" => rgb <= "100110";

when "010000101001001" => rgb <= "100110";

when "010000101001010" => rgb <= "100110";

when "010000101001011" => rgb <= "100110";

when "010000101001100" => rgb <= "100110";

when "010000101001101" => rgb <= "100110";

when "010000101001110" => rgb <= "100110";

when "010000101001111" => rgb <= "100110";

when "010000101010000" => rgb <= "100110";

when "010000101010001" => rgb <= "100110";

when "010000101010010" => rgb <= "100110";

when "010000101010011" => rgb <= "100110";

when "010000101010100" => rgb <= "100110";

when "010000101010101" => rgb <= "100110";

when "010000101010110" => rgb <= "100110";

when "010000101010111" => rgb <= "100110";

when "010000101011000" => rgb <= "100110";

when "010000101011001" => rgb <= "100110";

when "010000101011010" => rgb <= "100110";

when "010000101011011" => rgb <= "100110";

when "010000101011100" => rgb <= "100110";

when "010000101011101" => rgb <= "100110";

when "010000101011110" => rgb <= "100110";

when "010000101011111" => rgb <= "100110";

when "010000101100000" => rgb <= "100110";

when "010000101100001" => rgb <= "100110";

when "010000101100010" => rgb <= "100110";

when "010000101100011" => rgb <= "100110";

when "010000101100100" => rgb <= "100110";

when "010000101100101" => rgb <= "100110";

when "010000101100110" => rgb <= "100110";

when "010000101100111" => rgb <= "000000";

when "010001000111000" => rgb <= "000000";

when "010001000111001" => rgb <= "100110";

when "010001000111010" => rgb <= "100110";

when "010001000111011" => rgb <= "100110";

when "010001000111100" => rgb <= "100110";

when "010001000111101" => rgb <= "100110";

when "010001000111110" => rgb <= "100110";

when "010001000111111" => rgb <= "100110";

when "010001001000000" => rgb <= "100110";

when "010001001000001" => rgb <= "100110";

when "010001001000010" => rgb <= "100110";

when "010001001000011" => rgb <= "100110";

when "010001001000100" => rgb <= "100110";

when "010001001000101" => rgb <= "100110";

when "010001001000110" => rgb <= "100110";

when "010001001000111" => rgb <= "100110";

when "010001001001000" => rgb <= "100110";

when "010001001001001" => rgb <= "100110";

when "010001001001010" => rgb <= "100110";

when "010001001001011" => rgb <= "100110";

when "010001001001100" => rgb <= "100110";

when "010001001001101" => rgb <= "100110";

when "010001001001110" => rgb <= "100110";

when "010001001001111" => rgb <= "100110";

when "010001001010000" => rgb <= "100110";

when "010001001010001" => rgb <= "100110";

when "010001001010010" => rgb <= "100110";

when "010001001010011" => rgb <= "100110";

when "010001001010100" => rgb <= "100110";

when "010001001010101" => rgb <= "100110";

when "010001001010110" => rgb <= "100110";

when "010001001010111" => rgb <= "100110";

when "010001001011000" => rgb <= "100110";

when "010001001011001" => rgb <= "100110";

when "010001001011010" => rgb <= "100110";

when "010001001011011" => rgb <= "100110";

when "010001001011100" => rgb <= "100110";

when "010001001011101" => rgb <= "100110";

when "010001001011110" => rgb <= "100110";

when "010001001011111" => rgb <= "100110";

when "010001001100000" => rgb <= "100110";

when "010001001100001" => rgb <= "100110";

when "010001001100010" => rgb <= "100110";

when "010001001100011" => rgb <= "100110";

when "010001001100100" => rgb <= "100110";

when "010001001100101" => rgb <= "100110";

when "010001001100110" => rgb <= "100110";

when "010001001100111" => rgb <= "000000";

when "010001100111000" => rgb <= "000000";

when "010001100111001" => rgb <= "100110";

when "010001100111010" => rgb <= "100110";

when "010001100111011" => rgb <= "100110";

when "010001100111100" => rgb <= "100110";

when "010001100111101" => rgb <= "100110";

when "010001100111110" => rgb <= "100110";

when "010001100111111" => rgb <= "100110";

when "010001101000000" => rgb <= "100110";

when "010001101000001" => rgb <= "100110";

when "010001101000010" => rgb <= "100110";

when "010001101000011" => rgb <= "100110";

when "010001101000100" => rgb <= "100110";

when "010001101000101" => rgb <= "100110";

when "010001101000110" => rgb <= "100110";

when "010001101000111" => rgb <= "100110";

when "010001101001000" => rgb <= "100110";

when "010001101001001" => rgb <= "100110";

when "010001101001010" => rgb <= "100110";

when "010001101001011" => rgb <= "100110";

when "010001101001100" => rgb <= "100110";

when "010001101001101" => rgb <= "100110";

when "010001101001110" => rgb <= "100110";

when "010001101001111" => rgb <= "100110";

when "010001101010000" => rgb <= "100110";

when "010001101010001" => rgb <= "100110";

when "010001101010010" => rgb <= "100110";

when "010001101010011" => rgb <= "100110";

when "010001101010100" => rgb <= "100110";

when "010001101010101" => rgb <= "100110";

when "010001101010110" => rgb <= "100110";

when "010001101010111" => rgb <= "100110";

when "010001101011000" => rgb <= "100110";

when "010001101011001" => rgb <= "100110";

when "010001101011010" => rgb <= "100110";

when "010001101011011" => rgb <= "100110";

when "010001101011100" => rgb <= "100110";

when "010001101011101" => rgb <= "100110";

when "010001101011110" => rgb <= "100110";

when "010001101011111" => rgb <= "100110";

when "010001101100000" => rgb <= "100110";

when "010001101100001" => rgb <= "100110";

when "010001101100010" => rgb <= "100110";

when "010001101100011" => rgb <= "100110";

when "010001101100100" => rgb <= "100110";

when "010001101100101" => rgb <= "100110";

when "010001101100110" => rgb <= "100110";

when "010001101100111" => rgb <= "000000";

when "010010000111000" => rgb <= "000000";

when "010010000111001" => rgb <= "100110";

when "010010000111010" => rgb <= "100110";

when "010010000111011" => rgb <= "100110";

when "010010000111100" => rgb <= "100110";

when "010010000111101" => rgb <= "100110";

when "010010000111110" => rgb <= "100110";

when "010010000111111" => rgb <= "100110";

when "010010001000000" => rgb <= "100110";

when "010010001000001" => rgb <= "100110";

when "010010001000010" => rgb <= "100110";

when "010010001000011" => rgb <= "100110";

when "010010001000100" => rgb <= "100110";

when "010010001000101" => rgb <= "100110";

when "010010001000110" => rgb <= "100110";

when "010010001000111" => rgb <= "100110";

when "010010001001000" => rgb <= "100110";

when "010010001001001" => rgb <= "100110";

when "010010001001010" => rgb <= "100110";

when "010010001001011" => rgb <= "100110";

when "010010001001100" => rgb <= "100110";

when "010010001001101" => rgb <= "100110";

when "010010001001110" => rgb <= "100110";

when "010010001001111" => rgb <= "100110";

when "010010001010000" => rgb <= "100110";

when "010010001010001" => rgb <= "100110";

when "010010001010010" => rgb <= "100110";

when "010010001010011" => rgb <= "100110";

when "010010001010100" => rgb <= "100110";

when "010010001010101" => rgb <= "100110";

when "010010001010110" => rgb <= "100110";

when "010010001010111" => rgb <= "100110";

when "010010001011000" => rgb <= "100110";

when "010010001011001" => rgb <= "100110";

when "010010001011010" => rgb <= "100110";

when "010010001011011" => rgb <= "100110";

when "010010001011100" => rgb <= "100110";

when "010010001011101" => rgb <= "100110";

when "010010001011110" => rgb <= "100110";

when "010010001011111" => rgb <= "100110";

when "010010001100000" => rgb <= "100110";

when "010010001100001" => rgb <= "100110";

when "010010001100010" => rgb <= "100110";

when "010010001100011" => rgb <= "100110";

when "010010001100100" => rgb <= "100110";

when "010010001100101" => rgb <= "100110";

when "010010001100110" => rgb <= "100110";

when "010010001100111" => rgb <= "000000";

when "010010100111000" => rgb <= "000000";

when "010010100111001" => rgb <= "100110";

when "010010100111010" => rgb <= "100110";

when "010010100111011" => rgb <= "100110";

when "010010100111100" => rgb <= "100110";

when "010010100111101" => rgb <= "100110";

when "010010100111110" => rgb <= "100110";

when "010010100111111" => rgb <= "100110";

when "010010101000000" => rgb <= "100110";

when "010010101000001" => rgb <= "100110";

when "010010101000010" => rgb <= "100110";

when "010010101000011" => rgb <= "100110";

when "010010101000100" => rgb <= "100110";

when "010010101000101" => rgb <= "100110";

when "010010101000110" => rgb <= "100110";

when "010010101000111" => rgb <= "100110";

when "010010101001000" => rgb <= "100110";

when "010010101001001" => rgb <= "100110";

when "010010101001010" => rgb <= "100110";

when "010010101001011" => rgb <= "100110";

when "010010101001100" => rgb <= "100110";

when "010010101001101" => rgb <= "100110";

when "010010101001110" => rgb <= "100110";

when "010010101001111" => rgb <= "100110";

when "010010101010000" => rgb <= "100110";

when "010010101010001" => rgb <= "100110";

when "010010101010010" => rgb <= "100110";

when "010010101010011" => rgb <= "100110";

when "010010101010100" => rgb <= "100110";

when "010010101010101" => rgb <= "100110";

when "010010101010110" => rgb <= "100110";

when "010010101010111" => rgb <= "100110";

when "010010101011000" => rgb <= "100110";

when "010010101011001" => rgb <= "100110";

when "010010101011010" => rgb <= "100110";

when "010010101011011" => rgb <= "100110";

when "010010101011100" => rgb <= "100110";

when "010010101011101" => rgb <= "100110";

when "010010101011110" => rgb <= "100110";

when "010010101011111" => rgb <= "100110";

when "010010101100000" => rgb <= "100110";

when "010010101100001" => rgb <= "100110";

when "010010101100010" => rgb <= "100110";

when "010010101100011" => rgb <= "100110";

when "010010101100100" => rgb <= "100110";

when "010010101100101" => rgb <= "100110";

when "010010101100110" => rgb <= "100110";

when "010010101100111" => rgb <= "000000";

when "010011000111000" => rgb <= "000000";

when "010011000111001" => rgb <= "100110";

when "010011000111010" => rgb <= "100110";

when "010011000111011" => rgb <= "100110";

when "010011000111100" => rgb <= "100110";

when "010011000111101" => rgb <= "100110";

when "010011000111110" => rgb <= "100110";

when "010011000111111" => rgb <= "100110";

when "010011001000000" => rgb <= "000000";

when "010011001000001" => rgb <= "000000";

when "010011001000010" => rgb <= "000000";

when "010011001000011" => rgb <= "000000";

when "010011001000100" => rgb <= "000000";

when "010011001000101" => rgb <= "000000";

when "010011001000110" => rgb <= "000000";

when "010011001000111" => rgb <= "000000";

when "010011001001000" => rgb <= "000000";

when "010011001001001" => rgb <= "000000";

when "010011001001010" => rgb <= "000000";

when "010011001001011" => rgb <= "000000";

when "010011001001100" => rgb <= "000000";

when "010011001001101" => rgb <= "000000";

when "010011001001110" => rgb <= "000000";

when "010011001001111" => rgb <= "000000";

when "010011001010000" => rgb <= "000000";

when "010011001010001" => rgb <= "000000";

when "010011001010010" => rgb <= "000000";

when "010011001010011" => rgb <= "000000";

when "010011001010100" => rgb <= "000000";

when "010011001010101" => rgb <= "000000";

when "010011001010110" => rgb <= "000000";

when "010011001010111" => rgb <= "000000";

when "010011001011000" => rgb <= "000000";

when "010011001011001" => rgb <= "000000";

when "010011001011010" => rgb <= "000000";

when "010011001011011" => rgb <= "000000";

when "010011001011100" => rgb <= "000000";

when "010011001011101" => rgb <= "000000";

when "010011001011110" => rgb <= "000000";

when "010011001011111" => rgb <= "000000";

when "010011001100000" => rgb <= "000000";

when "010011001100001" => rgb <= "000000";

when "010011001100010" => rgb <= "000000";

when "010011001100011" => rgb <= "000000";

when "010011001100100" => rgb <= "000000";

when "010011001100101" => rgb <= "000000";

when "010011001100110" => rgb <= "000000";

when "010011001100111" => rgb <= "000000";

when "010011100111000" => rgb <= "000000";

when "010011100111001" => rgb <= "100110";

when "010011100111010" => rgb <= "100110";

when "010011100111011" => rgb <= "100110";

when "010011100111100" => rgb <= "100110";

when "010011100111101" => rgb <= "100110";

when "010011100111110" => rgb <= "100110";

when "010011100111111" => rgb <= "100110";

when "010011101000000" => rgb <= "000000";

when "010100000111000" => rgb <= "000000";

when "010100000111001" => rgb <= "100110";

when "010100000111010" => rgb <= "100110";

when "010100000111011" => rgb <= "100110";

when "010100000111100" => rgb <= "100110";

when "010100000111101" => rgb <= "100110";

when "010100000111110" => rgb <= "100110";

when "010100000111111" => rgb <= "100110";

when "010100001000000" => rgb <= "000000";

when "010100100111000" => rgb <= "000000";

when "010100100111001" => rgb <= "100110";

when "010100100111010" => rgb <= "100110";

when "010100100111011" => rgb <= "100110";

when "010100100111100" => rgb <= "100110";

when "010100100111101" => rgb <= "100110";

when "010100100111110" => rgb <= "100110";

when "010100100111111" => rgb <= "100110";

when "010100101000000" => rgb <= "000000";

when "010101000111000" => rgb <= "000000";

when "010101000111001" => rgb <= "100110";

when "010101000111010" => rgb <= "100110";

when "010101000111011" => rgb <= "100110";

when "010101000111100" => rgb <= "100110";

when "010101000111101" => rgb <= "100110";

when "010101000111110" => rgb <= "100110";

when "010101000111111" => rgb <= "100110";

when "010101001000000" => rgb <= "000000";

when "010101100111000" => rgb <= "000000";

when "010101100111001" => rgb <= "100110";

when "010101100111010" => rgb <= "100110";

when "010101100111011" => rgb <= "100110";

when "010101100111100" => rgb <= "100110";

when "010101100111101" => rgb <= "100110";

when "010101100111110" => rgb <= "100110";

when "010101100111111" => rgb <= "100110";

when "010101101000000" => rgb <= "000000";

when "010110000111000" => rgb <= "000000";

when "010110000111001" => rgb <= "100110";

when "010110000111010" => rgb <= "100110";

when "010110000111011" => rgb <= "100110";

when "010110000111100" => rgb <= "100110";

when "010110000111101" => rgb <= "100110";

when "010110000111110" => rgb <= "100110";

when "010110000111111" => rgb <= "100110";

when "010110001000000" => rgb <= "000000";

when "010110100111000" => rgb <= "000000";

when "010110100111001" => rgb <= "100110";

when "010110100111010" => rgb <= "100110";

when "010110100111011" => rgb <= "100110";

when "010110100111100" => rgb <= "100110";

when "010110100111101" => rgb <= "100110";

when "010110100111110" => rgb <= "100110";

when "010110100111111" => rgb <= "100110";

when "010110101000000" => rgb <= "000000";

when "010111000111000" => rgb <= "000000";

when "010111000111001" => rgb <= "100110";

when "010111000111010" => rgb <= "100110";

when "010111000111011" => rgb <= "100110";

when "010111000111100" => rgb <= "100110";

when "010111000111101" => rgb <= "100110";

when "010111000111110" => rgb <= "100110";

when "010111000111111" => rgb <= "100110";

when "010111001000000" => rgb <= "000000";

when "010111100111000" => rgb <= "000000";

when "010111100111001" => rgb <= "100110";

when "010111100111010" => rgb <= "100110";

when "010111100111011" => rgb <= "100110";

when "010111100111100" => rgb <= "100110";

when "010111100111101" => rgb <= "100110";

when "010111100111110" => rgb <= "100110";

when "010111100111111" => rgb <= "100110";

when "010111101000000" => rgb <= "000000";

when "011000000111000" => rgb <= "000000";

when "011000000111001" => rgb <= "100110";

when "011000000111010" => rgb <= "100110";

when "011000000111011" => rgb <= "100110";

when "011000000111100" => rgb <= "100110";

when "011000000111101" => rgb <= "100110";

when "011000000111110" => rgb <= "100110";

when "011000000111111" => rgb <= "100110";

when "011000001000000" => rgb <= "000000";

when "011000100111000" => rgb <= "000000";

when "011000100111001" => rgb <= "100110";

when "011000100111010" => rgb <= "100110";

when "011000100111011" => rgb <= "100110";

when "011000100111100" => rgb <= "100110";

when "011000100111101" => rgb <= "100110";

when "011000100111110" => rgb <= "100110";

when "011000100111111" => rgb <= "100110";

when "011000101000000" => rgb <= "000000";

when "011001000111000" => rgb <= "000000";

when "011001000111001" => rgb <= "100110";

when "011001000111010" => rgb <= "100110";

when "011001000111011" => rgb <= "100110";

when "011001000111100" => rgb <= "100110";

when "011001000111101" => rgb <= "100110";

when "011001000111110" => rgb <= "100110";

when "011001000111111" => rgb <= "100110";

when "011001001000000" => rgb <= "000000";

when "011001100111000" => rgb <= "000000";

when "011001100111001" => rgb <= "100110";

when "011001100111010" => rgb <= "100110";

when "011001100111011" => rgb <= "100110";

when "011001100111100" => rgb <= "100110";

when "011001100111101" => rgb <= "100110";

when "011001100111110" => rgb <= "100110";

when "011001100111111" => rgb <= "100110";

when "011001101000000" => rgb <= "000000";

when "011001101011111" => rgb <= "000000";

when "011001101100000" => rgb <= "000000";

when "011001101100001" => rgb <= "000000";

when "011001101100010" => rgb <= "000000";

when "011001101100011" => rgb <= "000000";

when "011001101100100" => rgb <= "000000";

when "011001101100101" => rgb <= "000000";

when "011001101100110" => rgb <= "000000";

when "011001101100111" => rgb <= "000000";

when "011010000111000" => rgb <= "000000";

when "011010000111001" => rgb <= "100110";

when "011010000111010" => rgb <= "100110";

when "011010000111011" => rgb <= "100110";

when "011010000111100" => rgb <= "100110";

when "011010000111101" => rgb <= "100110";

when "011010000111110" => rgb <= "100110";

when "011010000111111" => rgb <= "100110";

when "011010001000000" => rgb <= "000000";

when "011010001011111" => rgb <= "000000";

when "011010001100000" => rgb <= "100110";

when "011010001100001" => rgb <= "100110";

when "011010001100010" => rgb <= "100110";

when "011010001100011" => rgb <= "100110";

when "011010001100100" => rgb <= "100110";

when "011010001100101" => rgb <= "100110";

when "011010001100110" => rgb <= "100110";

when "011010001100111" => rgb <= "000000";

when "011010100111000" => rgb <= "000000";

when "011010100111001" => rgb <= "100110";

when "011010100111010" => rgb <= "100110";

when "011010100111011" => rgb <= "100110";

when "011010100111100" => rgb <= "100110";

when "011010100111101" => rgb <= "100110";

when "011010100111110" => rgb <= "100110";

when "011010100111111" => rgb <= "100110";

when "011010101000000" => rgb <= "000000";

when "011010101011111" => rgb <= "000000";

when "011010101100000" => rgb <= "100110";

when "011010101100001" => rgb <= "100110";

when "011010101100010" => rgb <= "100110";

when "011010101100011" => rgb <= "100110";

when "011010101100100" => rgb <= "100110";

when "011010101100101" => rgb <= "100110";

when "011010101100110" => rgb <= "100110";

when "011010101100111" => rgb <= "000000";

when "011011000111000" => rgb <= "000000";

when "011011000111001" => rgb <= "100110";

when "011011000111010" => rgb <= "100110";

when "011011000111011" => rgb <= "100110";

when "011011000111100" => rgb <= "100110";

when "011011000111101" => rgb <= "100110";

when "011011000111110" => rgb <= "100110";

when "011011000111111" => rgb <= "100110";

when "011011001000000" => rgb <= "000000";

when "011011001011111" => rgb <= "000000";

when "011011001100000" => rgb <= "100110";

when "011011001100001" => rgb <= "100110";

when "011011001100010" => rgb <= "100110";

when "011011001100011" => rgb <= "100110";

when "011011001100100" => rgb <= "100110";

when "011011001100101" => rgb <= "100110";

when "011011001100110" => rgb <= "100110";

when "011011001100111" => rgb <= "000000";

when "011011100111000" => rgb <= "000000";

when "011011100111001" => rgb <= "100110";

when "011011100111010" => rgb <= "100110";

when "011011100111011" => rgb <= "100110";

when "011011100111100" => rgb <= "100110";

when "011011100111101" => rgb <= "100110";

when "011011100111110" => rgb <= "100110";

when "011011100111111" => rgb <= "100110";

when "011011101000000" => rgb <= "000000";

when "011011101011111" => rgb <= "000000";

when "011011101100000" => rgb <= "100110";

when "011011101100001" => rgb <= "100110";

when "011011101100010" => rgb <= "100110";

when "011011101100011" => rgb <= "100110";

when "011011101100100" => rgb <= "100110";

when "011011101100101" => rgb <= "100110";

when "011011101100110" => rgb <= "100110";

when "011011101100111" => rgb <= "000000";

when "011100000111000" => rgb <= "000000";

when "011100000111001" => rgb <= "100110";

when "011100000111010" => rgb <= "100110";

when "011100000111011" => rgb <= "100110";

when "011100000111100" => rgb <= "100110";

when "011100000111101" => rgb <= "100110";

when "011100000111110" => rgb <= "100110";

when "011100000111111" => rgb <= "100110";

when "011100001000000" => rgb <= "000000";

when "011100001000001" => rgb <= "000000";

when "011100001000010" => rgb <= "000000";

when "011100001000011" => rgb <= "000000";

when "011100001000100" => rgb <= "000000";

when "011100001000101" => rgb <= "000000";

when "011100001000110" => rgb <= "000000";

when "011100001000111" => rgb <= "000000";

when "011100001001000" => rgb <= "000000";

when "011100001001001" => rgb <= "000000";

when "011100001001010" => rgb <= "000000";

when "011100001001011" => rgb <= "000000";

when "011100001001100" => rgb <= "000000";

when "011100001001101" => rgb <= "000000";

when "011100001001110" => rgb <= "000000";

when "011100001001111" => rgb <= "000000";

when "011100001010000" => rgb <= "000000";

when "011100001010001" => rgb <= "000000";

when "011100001010010" => rgb <= "000000";

when "011100001010011" => rgb <= "000000";

when "011100001010100" => rgb <= "000000";

when "011100001010101" => rgb <= "000000";

when "011100001010110" => rgb <= "000000";

when "011100001010111" => rgb <= "000000";

when "011100001011000" => rgb <= "000000";

when "011100001011001" => rgb <= "000000";

when "011100001011010" => rgb <= "000000";

when "011100001011011" => rgb <= "000000";

when "011100001011100" => rgb <= "000000";

when "011100001011101" => rgb <= "000000";

when "011100001011110" => rgb <= "000000";

when "011100001011111" => rgb <= "000000";

when "011100001100000" => rgb <= "100110";

when "011100001100001" => rgb <= "100110";

when "011100001100010" => rgb <= "100110";

when "011100001100011" => rgb <= "100110";

when "011100001100100" => rgb <= "100110";

when "011100001100101" => rgb <= "100110";

when "011100001100110" => rgb <= "100110";

when "011100001100111" => rgb <= "000000";

when "011100100111000" => rgb <= "000000";

when "011100100111001" => rgb <= "100110";

when "011100100111010" => rgb <= "100110";

when "011100100111011" => rgb <= "100110";

when "011100100111100" => rgb <= "100110";

when "011100100111101" => rgb <= "100110";

when "011100100111110" => rgb <= "100110";

when "011100100111111" => rgb <= "100110";

when "011100101000000" => rgb <= "100110";

when "011100101000001" => rgb <= "100110";

when "011100101000010" => rgb <= "100110";

when "011100101000011" => rgb <= "100110";

when "011100101000100" => rgb <= "100110";

when "011100101000101" => rgb <= "100110";

when "011100101000110" => rgb <= "100110";

when "011100101000111" => rgb <= "100110";

when "011100101001000" => rgb <= "100110";

when "011100101001001" => rgb <= "100110";

when "011100101001010" => rgb <= "100110";

when "011100101001011" => rgb <= "100110";

when "011100101001100" => rgb <= "100110";

when "011100101001101" => rgb <= "100110";

when "011100101001110" => rgb <= "100110";

when "011100101001111" => rgb <= "100110";

when "011100101010000" => rgb <= "100110";

when "011100101010001" => rgb <= "100110";

when "011100101010010" => rgb <= "100110";

when "011100101010011" => rgb <= "100110";

when "011100101010100" => rgb <= "100110";

when "011100101010101" => rgb <= "100110";

when "011100101010110" => rgb <= "100110";

when "011100101010111" => rgb <= "100110";

when "011100101011000" => rgb <= "100110";

when "011100101011001" => rgb <= "100110";

when "011100101011010" => rgb <= "100110";

when "011100101011011" => rgb <= "100110";

when "011100101011100" => rgb <= "100110";

when "011100101011101" => rgb <= "100110";

when "011100101011110" => rgb <= "100110";

when "011100101011111" => rgb <= "100110";

when "011100101100000" => rgb <= "100110";

when "011100101100001" => rgb <= "100110";

when "011100101100010" => rgb <= "100110";

when "011100101100011" => rgb <= "100110";

when "011100101100100" => rgb <= "100110";

when "011100101100101" => rgb <= "100110";

when "011100101100110" => rgb <= "100110";

when "011100101100111" => rgb <= "000000";

when "011101000111000" => rgb <= "000000";

when "011101000111001" => rgb <= "100110";

when "011101000111010" => rgb <= "100110";

when "011101000111011" => rgb <= "100110";

when "011101000111100" => rgb <= "100110";

when "011101000111101" => rgb <= "100110";

when "011101000111110" => rgb <= "100110";

when "011101000111111" => rgb <= "100110";

when "011101001000000" => rgb <= "100110";

when "011101001000001" => rgb <= "100110";

when "011101001000010" => rgb <= "100110";

when "011101001000011" => rgb <= "100110";

when "011101001000100" => rgb <= "100110";

when "011101001000101" => rgb <= "100110";

when "011101001000110" => rgb <= "100110";

when "011101001000111" => rgb <= "100110";

when "011101001001000" => rgb <= "100110";

when "011101001001001" => rgb <= "100110";

when "011101001001010" => rgb <= "100110";

when "011101001001011" => rgb <= "100110";

when "011101001001100" => rgb <= "100110";

when "011101001001101" => rgb <= "100110";

when "011101001001110" => rgb <= "100110";

when "011101001001111" => rgb <= "100110";

when "011101001010000" => rgb <= "100110";

when "011101001010001" => rgb <= "100110";

when "011101001010010" => rgb <= "100110";

when "011101001010011" => rgb <= "100110";

when "011101001010100" => rgb <= "100110";

when "011101001010101" => rgb <= "100110";

when "011101001010110" => rgb <= "100110";

when "011101001010111" => rgb <= "100110";

when "011101001011000" => rgb <= "100110";

when "011101001011001" => rgb <= "100110";

when "011101001011010" => rgb <= "100110";

when "011101001011011" => rgb <= "100110";

when "011101001011100" => rgb <= "100110";

when "011101001011101" => rgb <= "100110";

when "011101001011110" => rgb <= "100110";

when "011101001011111" => rgb <= "100110";

when "011101001100000" => rgb <= "100110";

when "011101001100001" => rgb <= "100110";

when "011101001100010" => rgb <= "100110";

when "011101001100011" => rgb <= "100110";

when "011101001100100" => rgb <= "100110";

when "011101001100101" => rgb <= "100110";

when "011101001100110" => rgb <= "100110";

when "011101001100111" => rgb <= "000000";

when "011101100111000" => rgb <= "000000";

when "011101100111001" => rgb <= "100110";

when "011101100111010" => rgb <= "100110";

when "011101100111011" => rgb <= "100110";

when "011101100111100" => rgb <= "100110";

when "011101100111101" => rgb <= "100110";

when "011101100111110" => rgb <= "100110";

when "011101100111111" => rgb <= "100110";

when "011101101000000" => rgb <= "100110";

when "011101101000001" => rgb <= "100110";

when "011101101000010" => rgb <= "100110";

when "011101101000011" => rgb <= "100110";

when "011101101000100" => rgb <= "100110";

when "011101101000101" => rgb <= "100110";

when "011101101000110" => rgb <= "100110";

when "011101101000111" => rgb <= "100110";

when "011101101001000" => rgb <= "100110";

when "011101101001001" => rgb <= "100110";

when "011101101001010" => rgb <= "100110";

when "011101101001011" => rgb <= "100110";

when "011101101001100" => rgb <= "100110";

when "011101101001101" => rgb <= "100110";

when "011101101001110" => rgb <= "100110";

when "011101101001111" => rgb <= "100110";

when "011101101010000" => rgb <= "100110";

when "011101101010001" => rgb <= "100110";

when "011101101010010" => rgb <= "100110";

when "011101101010011" => rgb <= "100110";

when "011101101010100" => rgb <= "100110";

when "011101101010101" => rgb <= "100110";

when "011101101010110" => rgb <= "100110";

when "011101101010111" => rgb <= "100110";

when "011101101011000" => rgb <= "100110";

when "011101101011001" => rgb <= "100110";

when "011101101011010" => rgb <= "100110";

when "011101101011011" => rgb <= "100110";

when "011101101011100" => rgb <= "100110";

when "011101101011101" => rgb <= "100110";

when "011101101011110" => rgb <= "100110";

when "011101101011111" => rgb <= "100110";

when "011101101100000" => rgb <= "100110";

when "011101101100001" => rgb <= "100110";

when "011101101100010" => rgb <= "100110";

when "011101101100011" => rgb <= "100110";

when "011101101100100" => rgb <= "100110";

when "011101101100101" => rgb <= "100110";

when "011101101100110" => rgb <= "100110";

when "011101101100111" => rgb <= "000000";

when "011110000111000" => rgb <= "000000";

when "011110000111001" => rgb <= "100110";

when "011110000111010" => rgb <= "100110";

when "011110000111011" => rgb <= "100110";

when "011110000111100" => rgb <= "100110";

when "011110000111101" => rgb <= "100110";

when "011110000111110" => rgb <= "100110";

when "011110000111111" => rgb <= "100110";

when "011110001000000" => rgb <= "100110";

when "011110001000001" => rgb <= "100110";

when "011110001000010" => rgb <= "100110";

when "011110001000011" => rgb <= "100110";

when "011110001000100" => rgb <= "100110";

when "011110001000101" => rgb <= "100110";

when "011110001000110" => rgb <= "100110";

when "011110001000111" => rgb <= "100110";

when "011110001001000" => rgb <= "100110";

when "011110001001001" => rgb <= "100110";

when "011110001001010" => rgb <= "100110";

when "011110001001011" => rgb <= "100110";

when "011110001001100" => rgb <= "100110";

when "011110001001101" => rgb <= "100110";

when "011110001001110" => rgb <= "100110";

when "011110001001111" => rgb <= "100110";

when "011110001010000" => rgb <= "100110";

when "011110001010001" => rgb <= "100110";

when "011110001010010" => rgb <= "100110";

when "011110001010011" => rgb <= "100110";

when "011110001010100" => rgb <= "100110";

when "011110001010101" => rgb <= "100110";

when "011110001010110" => rgb <= "100110";

when "011110001010111" => rgb <= "100110";

when "011110001011000" => rgb <= "100110";

when "011110001011001" => rgb <= "100110";

when "011110001011010" => rgb <= "100110";

when "011110001011011" => rgb <= "100110";

when "011110001011100" => rgb <= "100110";

when "011110001011101" => rgb <= "100110";

when "011110001011110" => rgb <= "100110";

when "011110001011111" => rgb <= "100110";

when "011110001100000" => rgb <= "100110";

when "011110001100001" => rgb <= "100110";

when "011110001100010" => rgb <= "100110";

when "011110001100011" => rgb <= "100110";

when "011110001100100" => rgb <= "100110";

when "011110001100101" => rgb <= "100110";

when "011110001100110" => rgb <= "100110";

when "011110001100111" => rgb <= "000000";

when "011110100111000" => rgb <= "000000";

when "011110100111001" => rgb <= "100110";

when "011110100111010" => rgb <= "100110";

when "011110100111011" => rgb <= "100110";

when "011110100111100" => rgb <= "100110";

when "011110100111101" => rgb <= "100110";

when "011110100111110" => rgb <= "100110";

when "011110100111111" => rgb <= "100110";

when "011110101000000" => rgb <= "100110";

when "011110101000001" => rgb <= "100110";

when "011110101000010" => rgb <= "100110";

when "011110101000011" => rgb <= "100110";

when "011110101000100" => rgb <= "100110";

when "011110101000101" => rgb <= "100110";

when "011110101000110" => rgb <= "100110";

when "011110101000111" => rgb <= "100110";

when "011110101001000" => rgb <= "100110";

when "011110101001001" => rgb <= "100110";

when "011110101001010" => rgb <= "100110";

when "011110101001011" => rgb <= "100110";

when "011110101001100" => rgb <= "100110";

when "011110101001101" => rgb <= "100110";

when "011110101001110" => rgb <= "100110";

when "011110101001111" => rgb <= "100110";

when "011110101010000" => rgb <= "100110";

when "011110101010001" => rgb <= "100110";

when "011110101010010" => rgb <= "100110";

when "011110101010011" => rgb <= "100110";

when "011110101010100" => rgb <= "100110";

when "011110101010101" => rgb <= "100110";

when "011110101010110" => rgb <= "100110";

when "011110101010111" => rgb <= "100110";

when "011110101011000" => rgb <= "100110";

when "011110101011001" => rgb <= "100110";

when "011110101011010" => rgb <= "100110";

when "011110101011011" => rgb <= "100110";

when "011110101011100" => rgb <= "100110";

when "011110101011101" => rgb <= "100110";

when "011110101011110" => rgb <= "100110";

when "011110101011111" => rgb <= "100110";

when "011110101100000" => rgb <= "100110";

when "011110101100001" => rgb <= "100110";

when "011110101100010" => rgb <= "100110";

when "011110101100011" => rgb <= "100110";

when "011110101100100" => rgb <= "100110";

when "011110101100101" => rgb <= "100110";

when "011110101100110" => rgb <= "100110";

when "011110101100111" => rgb <= "000000";

when "011111000111000" => rgb <= "000000";

when "011111000111001" => rgb <= "100110";

when "011111000111010" => rgb <= "100110";

when "011111000111011" => rgb <= "100110";

when "011111000111100" => rgb <= "100110";

when "011111000111101" => rgb <= "100110";

when "011111000111110" => rgb <= "100110";

when "011111000111111" => rgb <= "100110";

when "011111001000000" => rgb <= "100110";

when "011111001000001" => rgb <= "100110";

when "011111001000010" => rgb <= "100110";

when "011111001000011" => rgb <= "100110";

when "011111001000100" => rgb <= "100110";

when "011111001000101" => rgb <= "100110";

when "011111001000110" => rgb <= "100110";

when "011111001000111" => rgb <= "100110";

when "011111001001000" => rgb <= "100110";

when "011111001001001" => rgb <= "100110";

when "011111001001010" => rgb <= "100110";

when "011111001001011" => rgb <= "100110";

when "011111001001100" => rgb <= "100110";

when "011111001001101" => rgb <= "100110";

when "011111001001110" => rgb <= "100110";

when "011111001001111" => rgb <= "100110";

when "011111001010000" => rgb <= "100110";

when "011111001010001" => rgb <= "100110";

when "011111001010010" => rgb <= "100110";

when "011111001010011" => rgb <= "100110";

when "011111001010100" => rgb <= "100110";

when "011111001010101" => rgb <= "100110";

when "011111001010110" => rgb <= "100110";

when "011111001010111" => rgb <= "100110";

when "011111001011000" => rgb <= "100110";

when "011111001011001" => rgb <= "100110";

when "011111001011010" => rgb <= "100110";

when "011111001011011" => rgb <= "100110";

when "011111001011100" => rgb <= "100110";

when "011111001011101" => rgb <= "100110";

when "011111001011110" => rgb <= "100110";

when "011111001011111" => rgb <= "100110";

when "011111001100000" => rgb <= "100110";

when "011111001100001" => rgb <= "100110";

when "011111001100010" => rgb <= "100110";

when "011111001100011" => rgb <= "100110";

when "011111001100100" => rgb <= "100110";

when "011111001100101" => rgb <= "100110";

when "011111001100110" => rgb <= "100110";

when "011111001100111" => rgb <= "000000";

when "011111100111000" => rgb <= "000000";

when "011111100111001" => rgb <= "000000";

when "011111100111010" => rgb <= "000000";

when "011111100111011" => rgb <= "000000";

when "011111100111100" => rgb <= "000000";

when "011111100111101" => rgb <= "000000";

when "011111100111110" => rgb <= "000000";

when "011111100111111" => rgb <= "000000";

when "011111101000000" => rgb <= "000000";

when "011111101000001" => rgb <= "000000";

when "011111101000010" => rgb <= "000000";

when "011111101000011" => rgb <= "000000";

when "011111101000100" => rgb <= "000000";

when "011111101000101" => rgb <= "000000";

when "011111101000110" => rgb <= "000000";

when "011111101000111" => rgb <= "000000";

when "011111101001000" => rgb <= "000000";

when "011111101001001" => rgb <= "000000";

when "011111101001010" => rgb <= "000000";

when "011111101001011" => rgb <= "000000";

when "011111101001100" => rgb <= "000000";

when "011111101001101" => rgb <= "000000";

when "011111101001110" => rgb <= "000000";

when "011111101001111" => rgb <= "000000";

when "011111101010000" => rgb <= "000000";

when "011111101010001" => rgb <= "000000";

when "011111101010010" => rgb <= "000000";

when "011111101010011" => rgb <= "000000";

when "011111101010100" => rgb <= "000000";

when "011111101010101" => rgb <= "000000";

when "011111101010110" => rgb <= "000000";

when "011111101010111" => rgb <= "000000";

when "011111101011000" => rgb <= "000000";

when "011111101011001" => rgb <= "000000";

when "011111101011010" => rgb <= "000000";

when "011111101011011" => rgb <= "000000";

when "011111101011100" => rgb <= "000000";

when "011111101011101" => rgb <= "000000";

when "011111101011110" => rgb <= "000000";

when "011111101011111" => rgb <= "000000";

when "011111101100000" => rgb <= "000000";

when "011111101100001" => rgb <= "000000";

when "011111101100010" => rgb <= "000000";

when "011111101100011" => rgb <= "000000";

when "011111101100100" => rgb <= "000000";

when "011111101100101" => rgb <= "000000";

when "011111101100110" => rgb <= "000000";

when "011111101100111" => rgb <= "000000";
when others => rgb <= "111111"; --will update l8r
end case;
end if;
end process;
	addressOut <= address;
end;
