library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;


entity meow3 is --rom for the background
port(
    clk : in std_logic;
	address : in unsigned (14 downto 0); 
    rgb : out unsigned(5 downto 0)
);
end meow3;


architecture synth of meow3 is 

signal addressOut : unsigned(14 downto 0); 

begin
    process (clk) is begin
        if rising_edge(clk) then
            case addressOut is
                when "011010101011101" => rgb <= "000000";
		when "011010101011110" => rgb <= "000000";
		when "011010101011111" => rgb <= "000000";
		when "011010101100000" => rgb <= "000000";
		when "011010101100001" => rgb <= "000000";
		when "011010101100010" => rgb <= "000000";
		when "011010101100011" => rgb <= "000000";
		when "011010101100100" => rgb <= "000000";
		when "011010101100101" => rgb <= "000000";
		when "011010101100110" => rgb <= "000000";
		when "011010101100111" => rgb <= "000000";
		when "011010101101000" => rgb <= "000000";
		when "011010101101001" => rgb <= "000000";
		when "011010101101010" => rgb <= "000000";
		when "011010101101011" => rgb <= "000000";
		when "011010101101100" => rgb <= "000000";
		when "011010101101101" => rgb <= "000000";
		when "011010101101110" => rgb <= "000000";
		when "011010101101111" => rgb <= "000000";
		when "011010101110000" => rgb <= "000000";
		when "011010101110001" => rgb <= "000000";
		when "011010101110010" => rgb <= "000000";
		when "011010101110011" => rgb <= "000000";
		when "011011001011100" => rgb <= "000000";
		when "011011001011101" => rgb <= "111111";
		when "011011001011110" => rgb <= "111111";
		when "011011001011111" => rgb <= "111111";
		when "011011001100000" => rgb <= "111111";
		when "011011001100001" => rgb <= "111111";
		when "011011001100010" => rgb <= "111111";
		when "011011001100011" => rgb <= "111111";
		when "011011001100100" => rgb <= "111111";
		when "011011001100101" => rgb <= "111111";
		when "011011001100110" => rgb <= "111111";
		when "011011001100111" => rgb <= "111111";
		when "011011001101000" => rgb <= "111111";
		when "011011001101001" => rgb <= "111111";
		when "011011001101010" => rgb <= "111111";
		when "011011001101011" => rgb <= "111111";
		when "011011001101100" => rgb <= "111111";
		when "011011001101101" => rgb <= "111111";
		when "011011001101110" => rgb <= "111111";
		when "011011001101111" => rgb <= "111111";
		when "011011001110000" => rgb <= "111111";
		when "011011001110001" => rgb <= "111111";
		when "011011001110010" => rgb <= "111111";
		when "011011001110011" => rgb <= "111111";
		when "011011001110100" => rgb <= "000000";
		when "011011101011011" => rgb <= "000000";
		when "011011101011100" => rgb <= "111111";
		when "011011101011101" => rgb <= "111111";
		when "011011101011110" => rgb <= "111111";
		when "011011101011111" => rgb <= "111111";
		when "011011101100000" => rgb <= "111111";
		when "011011101100001" => rgb <= "111111";
		when "011011101100010" => rgb <= "111111";
		when "011011101100011" => rgb <= "111111";
		when "011011101100100" => rgb <= "111111";
		when "011011101100101" => rgb <= "111111";
		when "011011101100110" => rgb <= "111111";
		when "011011101100111" => rgb <= "111111";
		when "011011101101000" => rgb <= "111111";
		when "011011101101001" => rgb <= "111111";
		when "011011101101010" => rgb <= "111111";
		when "011011101101011" => rgb <= "111111";
		when "011011101101100" => rgb <= "111111";
		when "011011101101101" => rgb <= "111111";
		when "011011101101110" => rgb <= "111111";
		when "011011101101111" => rgb <= "111111";
		when "011011101110000" => rgb <= "111111";
		when "011011101110001" => rgb <= "111111";
		when "011011101110010" => rgb <= "111111";
		when "011011101110011" => rgb <= "111111";
		when "011011101110100" => rgb <= "111111";
		when "011011101110101" => rgb <= "000000";
		when "011100001011011" => rgb <= "000000";
		when "011100001011100" => rgb <= "111111";
		when "011100001011101" => rgb <= "111111";
		when "011100001011110" => rgb <= "111111";
		when "011100001011111" => rgb <= "000000";
		when "011100001100000" => rgb <= "000000";
		when "011100001100001" => rgb <= "000000";
		when "011100001100010" => rgb <= "000000";
		when "011100001100011" => rgb <= "111111";
		when "011100001100100" => rgb <= "111111";
		when "011100001100101" => rgb <= "000000";
		when "011100001100110" => rgb <= "000000";
		when "011100001100111" => rgb <= "000000";
		when "011100001101000" => rgb <= "111111";
		when "011100001101001" => rgb <= "000000";
		when "011100001101010" => rgb <= "000000";
		when "011100001101011" => rgb <= "000000";
		when "011100001101100" => rgb <= "111111";
		when "011100001101101" => rgb <= "000000";
		when "011100001101110" => rgb <= "111111";
		when "011100001101111" => rgb <= "111111";
		when "011100001110000" => rgb <= "111111";
		when "011100001110001" => rgb <= "000000";
		when "011100001110010" => rgb <= "111111";
		when "011100001110011" => rgb <= "111111";
		when "011100001110100" => rgb <= "111111";
		when "011100001110101" => rgb <= "000000";
		when "011100101011011" => rgb <= "000000";
		when "011100101011100" => rgb <= "111111";
		when "011100101011101" => rgb <= "111111";
		when "011100101011110" => rgb <= "111111";
		when "011100101011111" => rgb <= "000000";
		when "011100101100000" => rgb <= "111111";
		when "011100101100001" => rgb <= "000000";
		when "011100101100010" => rgb <= "111111";
		when "011100101100011" => rgb <= "000000";
		when "011100101100100" => rgb <= "111111";
		when "011100101100101" => rgb <= "000000";
		when "011100101100110" => rgb <= "111111";
		when "011100101100111" => rgb <= "111111";
		when "011100101101000" => rgb <= "111111";
		when "011100101101001" => rgb <= "000000";
		when "011100101101010" => rgb <= "111111";
		when "011100101101011" => rgb <= "000000";
		when "011100101101100" => rgb <= "111111";
		when "011100101101101" => rgb <= "000000";
		when "011100101101110" => rgb <= "111111";
		when "011100101101111" => rgb <= "111111";
		when "011100101110000" => rgb <= "111111";
		when "011100101110001" => rgb <= "000000";
		when "011100101110010" => rgb <= "111111";
		when "011100101110011" => rgb <= "111111";
		when "011100101110100" => rgb <= "111111";
		when "011100101110101" => rgb <= "000000";
		when "011101001011011" => rgb <= "000000";
		when "011101001011100" => rgb <= "111111";
		when "011101001011101" => rgb <= "111111";
		when "011101001011110" => rgb <= "111111";
		when "011101001011111" => rgb <= "000000";
		when "011101001100000" => rgb <= "111111";
		when "011101001100001" => rgb <= "000000";
		when "011101001100010" => rgb <= "111111";
		when "011101001100011" => rgb <= "000000";
		when "011101001100100" => rgb <= "111111";
		when "011101001100101" => rgb <= "000000";
		when "011101001100110" => rgb <= "000000";
		when "011101001100111" => rgb <= "111111";
		when "011101001101000" => rgb <= "111111";
		when "011101001101001" => rgb <= "000000";
		when "011101001101010" => rgb <= "111111";
		when "011101001101011" => rgb <= "000000";
		when "011101001101100" => rgb <= "111111";
		when "011101001101101" => rgb <= "000000";
		when "011101001101110" => rgb <= "111111";
		when "011101001101111" => rgb <= "000000";
		when "011101001110000" => rgb <= "111111";
		when "011101001110001" => rgb <= "000000";
		when "011101001110010" => rgb <= "111111";
		when "011101001110011" => rgb <= "111111";
		when "011101001110100" => rgb <= "111111";
		when "011101001110101" => rgb <= "000000";
		when "011101101011011" => rgb <= "000000";
		when "011101101011100" => rgb <= "111111";
		when "011101101011101" => rgb <= "111111";
		when "011101101011110" => rgb <= "111111";
		when "011101101011111" => rgb <= "000000";
		when "011101101100000" => rgb <= "111111";
		when "011101101100001" => rgb <= "000000";
		when "011101101100010" => rgb <= "111111";
		when "011101101100011" => rgb <= "000000";
		when "011101101100100" => rgb <= "111111";
		when "011101101100101" => rgb <= "000000";
		when "011101101100110" => rgb <= "111111";
		when "011101101100111" => rgb <= "111111";
		when "011101101101000" => rgb <= "111111";
		when "011101101101001" => rgb <= "000000";
		when "011101101101010" => rgb <= "111111";
		when "011101101101011" => rgb <= "000000";
		when "011101101101100" => rgb <= "111111";
		when "011101101101101" => rgb <= "000000";
		when "011101101101110" => rgb <= "111111";
		when "011101101101111" => rgb <= "000000";
		when "011101101110000" => rgb <= "111111";
		when "011101101110001" => rgb <= "000000";
		when "011101101110010" => rgb <= "111111";
		when "011101101110011" => rgb <= "111111";
		when "011101101110100" => rgb <= "111111";
		when "011101101110101" => rgb <= "000000";
		when "011110001011011" => rgb <= "000000";
		when "011110001011100" => rgb <= "111111";
		when "011110001011101" => rgb <= "111111";
		when "011110001011110" => rgb <= "111111";
		when "011110001011111" => rgb <= "000000";
		when "011110001100000" => rgb <= "111111";
		when "011110001100001" => rgb <= "000000";
		when "011110001100010" => rgb <= "111111";
		when "011110001100011" => rgb <= "000000";
		when "011110001100100" => rgb <= "111111";
		when "011110001100101" => rgb <= "000000";
		when "011110001100110" => rgb <= "000000";
		when "011110001100111" => rgb <= "000000";
		when "011110001101000" => rgb <= "111111";
		when "011110001101001" => rgb <= "000000";
		when "011110001101010" => rgb <= "000000";
		when "011110001101011" => rgb <= "000000";
		when "011110001101100" => rgb <= "111111";
		when "011110001101101" => rgb <= "000000";
		when "011110001101110" => rgb <= "000000";
		when "011110001101111" => rgb <= "000000";
		when "011110001110000" => rgb <= "000000";
		when "011110001110001" => rgb <= "111111";
		when "011110001110010" => rgb <= "111111";
		when "011110001110011" => rgb <= "111111";
		when "011110001110100" => rgb <= "111111";
		when "011110001110101" => rgb <= "000000";
		when "011110101011011" => rgb <= "000000";
		when "011110101011100" => rgb <= "000000";
		when "011110101011101" => rgb <= "111111";
		when "011110101011110" => rgb <= "111111";
		when "011110101011111" => rgb <= "111111";
		when "011110101100000" => rgb <= "111111";
		when "011110101100001" => rgb <= "111111";
		when "011110101100010" => rgb <= "111111";
		when "011110101100011" => rgb <= "111111";
		when "011110101100100" => rgb <= "111111";
		when "011110101100101" => rgb <= "111111";
		when "011110101100110" => rgb <= "111111";
		when "011110101100111" => rgb <= "111111";
		when "011110101101000" => rgb <= "111111";
		when "011110101101001" => rgb <= "111111";
		when "011110101101010" => rgb <= "111111";
		when "011110101101011" => rgb <= "111111";
		when "011110101101100" => rgb <= "111111";
		when "011110101101101" => rgb <= "111111";
		when "011110101101110" => rgb <= "111111";
		when "011110101101111" => rgb <= "111111";
		when "011110101110000" => rgb <= "111111";
		when "011110101110001" => rgb <= "111111";
		when "011110101110010" => rgb <= "111111";
		when "011110101110011" => rgb <= "111111";
		when "011110101110100" => rgb <= "111111";
		when "011110101110101" => rgb <= "000000";
		when "011111001011100" => rgb <= "000000";
		when "011111001011101" => rgb <= "111111";
		when "011111001011110" => rgb <= "111111";
		when "011111001011111" => rgb <= "111111";
		when "011111001100000" => rgb <= "111111";
		when "011111001100001" => rgb <= "111111";
		when "011111001100010" => rgb <= "111111";
		when "011111001100011" => rgb <= "111111";
		when "011111001100100" => rgb <= "111111";
		when "011111001100101" => rgb <= "111111";
		when "011111001100110" => rgb <= "111111";
		when "011111001100111" => rgb <= "111111";
		when "011111001101000" => rgb <= "111111";
		when "011111001101001" => rgb <= "111111";
		when "011111001101010" => rgb <= "111111";
		when "011111001101011" => rgb <= "111111";
		when "011111001101100" => rgb <= "111111";
		when "011111001101101" => rgb <= "111111";
		when "011111001101110" => rgb <= "111111";
		when "011111001101111" => rgb <= "111111";
		when "011111001110000" => rgb <= "111111";
		when "011111001110001" => rgb <= "111111";
		when "011111001110010" => rgb <= "111111";
		when "011111001110011" => rgb <= "111111";
		when "011111001110100" => rgb <= "000000";
		when "011111101011101" => rgb <= "000000";
		when "011111101011110" => rgb <= "000000";
		when "011111101011111" => rgb <= "000000";
		when "011111101100000" => rgb <= "000000";
		when "011111101100001" => rgb <= "111111";
		when "011111101100010" => rgb <= "111111";
		when "011111101100011" => rgb <= "111111";
		when "011111101100100" => rgb <= "000000";
		when "011111101100101" => rgb <= "000000";
		when "011111101100110" => rgb <= "000000";
		when "011111101100111" => rgb <= "000000";
		when "011111101101000" => rgb <= "000000";
		when "011111101101001" => rgb <= "000000";
		when "011111101101010" => rgb <= "000000";
		when "011111101101011" => rgb <= "000000";
		when "011111101101100" => rgb <= "000000";
		when "011111101101101" => rgb <= "000000";
		when "011111101101110" => rgb <= "000000";
		when "011111101101111" => rgb <= "000000";
		when "011111101110000" => rgb <= "000000";
		when "011111101110001" => rgb <= "000000";
		when "011111101110010" => rgb <= "000000";
		when "011111101110011" => rgb <= "000000";
		when "100000001100000" => rgb <= "000000";
		when "100000001100001" => rgb <= "111111";
		when "100000001100010" => rgb <= "111111";
		when "100000001100011" => rgb <= "111111";
		when "100000001100100" => rgb <= "000000";
		when "100000101011111" => rgb <= "000000";
		when "100000101100000" => rgb <= "111111";
		when "100000101100001" => rgb <= "111111";
		when "100000101100010" => rgb <= "111111";
		when "100000101100011" => rgb <= "000000";
		when "100001001011111" => rgb <= "000000";
		when "100001001100000" => rgb <= "111111";
		when "100001001100001" => rgb <= "111111";
		when "100001001100010" => rgb <= "000000";
		when "100001101011111" => rgb <= "000000";
		when "100001101100000" => rgb <= "000000";
		when "100001101100001" => rgb <= "000000";
		when others => rgb <= "110000";
	end case;
end if;
end process;
	addressOut <= address;
end; 
