library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;


entity yourturn is 
port(
    clk : in std_logic;
	address : in unsigned (14 downto 0); 
    rgb : out unsigned(5 downto 0)
);
end yourturn;


architecture synth of yourturn is 

signal addressOut : unsigned(14 downto 0); 

begin
    process (clk) is begin
        if rising_edge(clk) then
            case addressOut is
			when "001001000101101" => rgb <= "000000";

when "001001000101110" => rgb <= "000000";

when "001001000101111" => rgb <= "000000";

when "001001000110000" => rgb <= "000000";

when "001001000110001" => rgb <= "000000";

when "001001000110110" => rgb <= "000000";

when "001001000110111" => rgb <= "000000";

when "001001000111000" => rgb <= "000000";

when "001001000111001" => rgb <= "000000";

when "001001000111010" => rgb <= "000000";

when "001001001000000" => rgb <= "000000";

when "001001001000001" => rgb <= "000000";

when "001001001000010" => rgb <= "000000";

when "001001001000011" => rgb <= "000000";

when "001001001000100" => rgb <= "000000";

when "001001001000101" => rgb <= "000000";

when "001001001000110" => rgb <= "000000";

when "001001001000111" => rgb <= "000000";

when "001001001001101" => rgb <= "000000";

when "001001001001110" => rgb <= "000000";

when "001001001001111" => rgb <= "000000";

when "001001001010000" => rgb <= "000000";

when "001001001010001" => rgb <= "000000";

when "001001001010110" => rgb <= "000000";

when "001001001010111" => rgb <= "000000";

when "001001001011000" => rgb <= "000000";

when "001001001011001" => rgb <= "000000";

when "001001001011010" => rgb <= "000000";

when "001001001011101" => rgb <= "000000";

when "001001001011110" => rgb <= "000000";

when "001001001011111" => rgb <= "000000";

when "001001001100000" => rgb <= "000000";

when "001001001100001" => rgb <= "000000";

when "001001001100010" => rgb <= "000000";

when "001001001100011" => rgb <= "000000";

when "001001001100100" => rgb <= "000000";

when "001001001100101" => rgb <= "000000";

when "001001001100110" => rgb <= "000000";

when "001001001100111" => rgb <= "000000";

when "001001100101101" => rgb <= "000000";

when "001001100101110" => rgb <= "100110";

when "001001100101111" => rgb <= "100110";

when "001001100110000" => rgb <= "100110";

when "001001100110001" => rgb <= "000000";

when "001001100110110" => rgb <= "000000";

when "001001100110111" => rgb <= "100110";

when "001001100111000" => rgb <= "100110";

when "001001100111001" => rgb <= "100110";

when "001001100111010" => rgb <= "000000";

when "001001100111110" => rgb <= "000000";

when "001001100111111" => rgb <= "000000";

when "001001101000000" => rgb <= "000000";

when "001001101000001" => rgb <= "100110";

when "001001101000010" => rgb <= "100110";

when "001001101000011" => rgb <= "100110";

when "001001101000100" => rgb <= "100110";

when "001001101000101" => rgb <= "100110";

when "001001101000110" => rgb <= "100110";

when "001001101000111" => rgb <= "000000";

when "001001101001000" => rgb <= "000000";

when "001001101001001" => rgb <= "000000";

when "001001101001101" => rgb <= "000000";

when "001001101001110" => rgb <= "100110";

when "001001101001111" => rgb <= "100110";

when "001001101010000" => rgb <= "100110";

when "001001101010001" => rgb <= "000000";

when "001001101010110" => rgb <= "000000";

when "001001101010111" => rgb <= "100110";

when "001001101011000" => rgb <= "100110";

when "001001101011001" => rgb <= "100110";

when "001001101011010" => rgb <= "000000";

when "001001101011101" => rgb <= "000000";

when "001001101011110" => rgb <= "100110";

when "001001101011111" => rgb <= "100110";

when "001001101100000" => rgb <= "100110";

when "001001101100001" => rgb <= "100110";

when "001001101100010" => rgb <= "100110";

when "001001101100011" => rgb <= "100110";

when "001001101100100" => rgb <= "100110";

when "001001101100101" => rgb <= "100110";

when "001001101100110" => rgb <= "100110";

when "001001101100111" => rgb <= "000000";

when "001001101101000" => rgb <= "000000";

when "001001101101001" => rgb <= "000000";

when "001010000101101" => rgb <= "000000";

when "001010000101110" => rgb <= "100110";

when "001010000101111" => rgb <= "100110";

when "001010000110000" => rgb <= "100110";

when "001010000110001" => rgb <= "000000";

when "001010000110110" => rgb <= "000000";

when "001010000110111" => rgb <= "100110";

when "001010000111000" => rgb <= "100110";

when "001010000111001" => rgb <= "100110";

when "001010000111010" => rgb <= "000000";

when "001010000111110" => rgb <= "000000";

when "001010000111111" => rgb <= "100110";

when "001010001000000" => rgb <= "100110";

when "001010001000001" => rgb <= "100110";

when "001010001000010" => rgb <= "100110";

when "001010001000011" => rgb <= "100110";

when "001010001000100" => rgb <= "100110";

when "001010001000101" => rgb <= "100110";

when "001010001000110" => rgb <= "100110";

when "001010001000111" => rgb <= "100110";

when "001010001001000" => rgb <= "100110";

when "001010001001001" => rgb <= "000000";

when "001010001001101" => rgb <= "000000";

when "001010001001110" => rgb <= "100110";

when "001010001001111" => rgb <= "100110";

when "001010001010000" => rgb <= "100110";

when "001010001010001" => rgb <= "000000";

when "001010001010110" => rgb <= "000000";

when "001010001010111" => rgb <= "100110";

when "001010001011000" => rgb <= "100110";

when "001010001011001" => rgb <= "100110";

when "001010001011010" => rgb <= "000000";

when "001010001011101" => rgb <= "000000";

when "001010001011110" => rgb <= "100110";

when "001010001011111" => rgb <= "100110";

when "001010001100000" => rgb <= "100110";

when "001010001100001" => rgb <= "100110";

when "001010001100010" => rgb <= "100110";

when "001010001100011" => rgb <= "100110";

when "001010001100100" => rgb <= "100110";

when "001010001100101" => rgb <= "100110";

when "001010001100110" => rgb <= "100110";

when "001010001100111" => rgb <= "100110";

when "001010001101000" => rgb <= "100110";

when "001010001101001" => rgb <= "000000";

when "001010100101101" => rgb <= "000000";

when "001010100101110" => rgb <= "100110";

when "001010100101111" => rgb <= "100110";

when "001010100110000" => rgb <= "100110";

when "001010100110001" => rgb <= "000000";

when "001010100110110" => rgb <= "000000";

when "001010100110111" => rgb <= "100110";

when "001010100111000" => rgb <= "100110";

when "001010100111001" => rgb <= "100110";

when "001010100111010" => rgb <= "000000";

when "001010100111101" => rgb <= "000000";

when "001010100111110" => rgb <= "000000";

when "001010100111111" => rgb <= "100110";

when "001010101000000" => rgb <= "100110";

when "001010101000001" => rgb <= "100110";

when "001010101000010" => rgb <= "100110";

when "001010101000011" => rgb <= "100110";

when "001010101000100" => rgb <= "100110";

when "001010101000101" => rgb <= "100110";

when "001010101000110" => rgb <= "100110";

when "001010101000111" => rgb <= "100110";

when "001010101001000" => rgb <= "100110";

when "001010101001001" => rgb <= "000000";

when "001010101001010" => rgb <= "000000";

when "001010101001101" => rgb <= "000000";

when "001010101001110" => rgb <= "100110";

when "001010101001111" => rgb <= "100110";

when "001010101010000" => rgb <= "100110";

when "001010101010001" => rgb <= "000000";

when "001010101010110" => rgb <= "000000";

when "001010101010111" => rgb <= "100110";

when "001010101011000" => rgb <= "100110";

when "001010101011001" => rgb <= "100110";

when "001010101011010" => rgb <= "000000";

when "001010101011101" => rgb <= "000000";

when "001010101011110" => rgb <= "100110";

when "001010101011111" => rgb <= "100110";

when "001010101100000" => rgb <= "100110";

when "001010101100001" => rgb <= "000000";

when "001010101100010" => rgb <= "000000";

when "001010101100011" => rgb <= "000000";

when "001010101100100" => rgb <= "000000";

when "001010101100101" => rgb <= "000000";

when "001010101100110" => rgb <= "100110";

when "001010101100111" => rgb <= "100110";

when "001010101101000" => rgb <= "100110";

when "001010101101001" => rgb <= "000000";

when "001011000101101" => rgb <= "000000";

when "001011000101110" => rgb <= "100110";

when "001011000101111" => rgb <= "100110";

when "001011000110000" => rgb <= "100110";

when "001011000110001" => rgb <= "000000";

when "001011000110010" => rgb <= "000000";

when "001011000110101" => rgb <= "000000";

when "001011000110110" => rgb <= "000000";

when "001011000110111" => rgb <= "100110";

when "001011000111000" => rgb <= "100110";

when "001011000111001" => rgb <= "100110";

when "001011000111010" => rgb <= "000000";

when "001011000111101" => rgb <= "000000";

when "001011000111110" => rgb <= "100110";

when "001011000111111" => rgb <= "100110";

when "001011001000000" => rgb <= "100110";

when "001011001000001" => rgb <= "100110";

when "001011001000010" => rgb <= "000000";

when "001011001000011" => rgb <= "000000";

when "001011001000100" => rgb <= "000000";

when "001011001000101" => rgb <= "000000";

when "001011001000110" => rgb <= "100110";

when "001011001000111" => rgb <= "100110";

when "001011001001000" => rgb <= "100110";

when "001011001001001" => rgb <= "100110";

when "001011001001010" => rgb <= "000000";

when "001011001001101" => rgb <= "000000";

when "001011001001110" => rgb <= "100110";

when "001011001001111" => rgb <= "100110";

when "001011001010000" => rgb <= "100110";

when "001011001010001" => rgb <= "000000";

when "001011001010110" => rgb <= "000000";

when "001011001010111" => rgb <= "100110";

when "001011001011000" => rgb <= "100110";

when "001011001011001" => rgb <= "100110";

when "001011001011010" => rgb <= "000000";

when "001011001011101" => rgb <= "000000";

when "001011001011110" => rgb <= "100110";

when "001011001011111" => rgb <= "100110";

when "001011001100000" => rgb <= "100110";

when "001011001100001" => rgb <= "000000";

when "001011001100101" => rgb <= "000000";

when "001011001100110" => rgb <= "100110";

when "001011001100111" => rgb <= "100110";

when "001011001101000" => rgb <= "100110";

when "001011001101001" => rgb <= "000000";

when "001011100101101" => rgb <= "000000";

when "001011100101110" => rgb <= "100110";

when "001011100101111" => rgb <= "100110";

when "001011100110000" => rgb <= "100110";

when "001011100110001" => rgb <= "100110";

when "001011100110010" => rgb <= "000000";

when "001011100110101" => rgb <= "000000";

when "001011100110110" => rgb <= "100110";

when "001011100110111" => rgb <= "100110";

when "001011100111000" => rgb <= "100110";

when "001011100111001" => rgb <= "100110";

when "001011100111010" => rgb <= "000000";

when "001011100111101" => rgb <= "000000";

when "001011100111110" => rgb <= "100110";

when "001011100111111" => rgb <= "100110";

when "001011101000000" => rgb <= "100110";

when "001011101000001" => rgb <= "000000";

when "001011101000010" => rgb <= "000000";

when "001011101000101" => rgb <= "000000";

when "001011101000110" => rgb <= "000000";

when "001011101000111" => rgb <= "100110";

when "001011101001000" => rgb <= "100110";

when "001011101001001" => rgb <= "100110";

when "001011101001010" => rgb <= "000000";

when "001011101001101" => rgb <= "000000";

when "001011101001110" => rgb <= "100110";

when "001011101001111" => rgb <= "100110";

when "001011101010000" => rgb <= "100110";

when "001011101010001" => rgb <= "000000";

when "001011101010110" => rgb <= "000000";

when "001011101010111" => rgb <= "100110";

when "001011101011000" => rgb <= "100110";

when "001011101011001" => rgb <= "100110";

when "001011101011010" => rgb <= "000000";

when "001011101011101" => rgb <= "000000";

when "001011101011110" => rgb <= "100110";

when "001011101011111" => rgb <= "100110";

when "001011101100000" => rgb <= "100110";

when "001011101100001" => rgb <= "000000";

when "001011101100101" => rgb <= "000000";

when "001011101100110" => rgb <= "100110";

when "001011101100111" => rgb <= "100110";

when "001011101101000" => rgb <= "100110";

when "001011101101001" => rgb <= "000000";

when "001100000101101" => rgb <= "000000";

when "001100000101110" => rgb <= "000000";

when "001100000101111" => rgb <= "100110";

when "001100000110000" => rgb <= "100110";

when "001100000110001" => rgb <= "100110";

when "001100000110010" => rgb <= "000000";

when "001100000110011" => rgb <= "000000";

when "001100000110100" => rgb <= "000000";

when "001100000110101" => rgb <= "000000";

when "001100000110110" => rgb <= "100110";

when "001100000110111" => rgb <= "100110";

when "001100000111000" => rgb <= "100110";

when "001100000111001" => rgb <= "000000";

when "001100000111010" => rgb <= "000000";

when "001100000111101" => rgb <= "000000";

when "001100000111110" => rgb <= "100110";

when "001100000111111" => rgb <= "100110";

when "001100001000000" => rgb <= "100110";

when "001100001000001" => rgb <= "000000";

when "001100001000110" => rgb <= "000000";

when "001100001000111" => rgb <= "100110";

when "001100001001000" => rgb <= "100110";

when "001100001001001" => rgb <= "100110";

when "001100001001010" => rgb <= "000000";

when "001100001001101" => rgb <= "000000";

when "001100001001110" => rgb <= "100110";

when "001100001001111" => rgb <= "100110";

when "001100001010000" => rgb <= "100110";

when "001100001010001" => rgb <= "000000";

when "001100001010110" => rgb <= "000000";

when "001100001010111" => rgb <= "100110";

when "001100001011000" => rgb <= "100110";

when "001100001011001" => rgb <= "100110";

when "001100001011010" => rgb <= "000000";

when "001100001011101" => rgb <= "000000";

when "001100001011110" => rgb <= "100110";

when "001100001011111" => rgb <= "100110";

when "001100001100000" => rgb <= "100110";

when "001100001100001" => rgb <= "000000";

when "001100001100100" => rgb <= "000000";

when "001100001100101" => rgb <= "000000";

when "001100001100110" => rgb <= "100110";

when "001100001100111" => rgb <= "100110";

when "001100001101000" => rgb <= "100110";

when "001100001101001" => rgb <= "000000";

when "001100100101110" => rgb <= "000000";

when "001100100101111" => rgb <= "100110";

when "001100100110000" => rgb <= "100110";

when "001100100110001" => rgb <= "100110";

when "001100100110010" => rgb <= "100110";

when "001100100110011" => rgb <= "100110";

when "001100100110100" => rgb <= "100110";

when "001100100110101" => rgb <= "100110";

when "001100100110110" => rgb <= "100110";

when "001100100110111" => rgb <= "100110";

when "001100100111000" => rgb <= "100110";

when "001100100111001" => rgb <= "000000";

when "001100100111101" => rgb <= "000000";

when "001100100111110" => rgb <= "100110";

when "001100100111111" => rgb <= "100110";

when "001100101000000" => rgb <= "100110";

when "001100101000001" => rgb <= "000000";

when "001100101000110" => rgb <= "000000";

when "001100101000111" => rgb <= "100110";

when "001100101001000" => rgb <= "100110";

when "001100101001001" => rgb <= "100110";

when "001100101001010" => rgb <= "000000";

when "001100101001101" => rgb <= "000000";

when "001100101001110" => rgb <= "100110";

when "001100101001111" => rgb <= "100110";

when "001100101010000" => rgb <= "100110";

when "001100101010001" => rgb <= "000000";

when "001100101010110" => rgb <= "000000";

when "001100101010111" => rgb <= "100110";

when "001100101011000" => rgb <= "100110";

when "001100101011001" => rgb <= "100110";

when "001100101011010" => rgb <= "000000";

when "001100101011101" => rgb <= "000000";

when "001100101011110" => rgb <= "100110";

when "001100101011111" => rgb <= "100110";

when "001100101100000" => rgb <= "100110";

when "001100101100001" => rgb <= "000000";

when "001100101100010" => rgb <= "000000";

when "001100101100011" => rgb <= "000000";

when "001100101100100" => rgb <= "000000";

when "001100101100101" => rgb <= "100110";

when "001100101100110" => rgb <= "100110";

when "001100101100111" => rgb <= "100110";

when "001100101101000" => rgb <= "100110";

when "001100101101001" => rgb <= "000000";

when "001101000101110" => rgb <= "000000";

when "001101000101111" => rgb <= "000000";

when "001101000110000" => rgb <= "100110";

when "001101000110001" => rgb <= "100110";

when "001101000110010" => rgb <= "100110";

when "001101000110011" => rgb <= "100110";

when "001101000110100" => rgb <= "100110";

when "001101000110101" => rgb <= "100110";

when "001101000110110" => rgb <= "100110";

when "001101000110111" => rgb <= "100110";

when "001101000111000" => rgb <= "000000";

when "001101000111001" => rgb <= "000000";

when "001101000111101" => rgb <= "000000";

when "001101000111110" => rgb <= "100110";

when "001101000111111" => rgb <= "100110";

when "001101001000000" => rgb <= "100110";

when "001101001000001" => rgb <= "000000";

when "001101001000110" => rgb <= "000000";

when "001101001000111" => rgb <= "100110";

when "001101001001000" => rgb <= "100110";

when "001101001001001" => rgb <= "100110";

when "001101001001010" => rgb <= "000000";

when "001101001001101" => rgb <= "000000";

when "001101001001110" => rgb <= "100110";

when "001101001001111" => rgb <= "100110";

when "001101001010000" => rgb <= "100110";

when "001101001010001" => rgb <= "000000";

when "001101001010110" => rgb <= "000000";

when "001101001010111" => rgb <= "100110";

when "001101001011000" => rgb <= "100110";

when "001101001011001" => rgb <= "100110";

when "001101001011010" => rgb <= "000000";

when "001101001011101" => rgb <= "000000";

when "001101001011110" => rgb <= "100110";

when "001101001011111" => rgb <= "100110";

when "001101001100000" => rgb <= "100110";

when "001101001100001" => rgb <= "100110";

when "001101001100010" => rgb <= "100110";

when "001101001100011" => rgb <= "100110";

when "001101001100100" => rgb <= "100110";

when "001101001100101" => rgb <= "100110";

when "001101001100110" => rgb <= "100110";

when "001101001100111" => rgb <= "000000";

when "001101001101000" => rgb <= "000000";

when "001101001101001" => rgb <= "000000";

when "001101100101111" => rgb <= "000000";

when "001101100110000" => rgb <= "000000";

when "001101100110001" => rgb <= "000000";

when "001101100110010" => rgb <= "100110";

when "001101100110011" => rgb <= "100110";

when "001101100110100" => rgb <= "100110";

when "001101100110101" => rgb <= "100110";

when "001101100110110" => rgb <= "000000";

when "001101100110111" => rgb <= "000000";

when "001101100111000" => rgb <= "000000";

when "001101100111101" => rgb <= "000000";

when "001101100111110" => rgb <= "100110";

when "001101100111111" => rgb <= "100110";

when "001101101000000" => rgb <= "100110";

when "001101101000001" => rgb <= "000000";

when "001101101000110" => rgb <= "000000";

when "001101101000111" => rgb <= "100110";

when "001101101001000" => rgb <= "100110";

when "001101101001001" => rgb <= "100110";

when "001101101001010" => rgb <= "000000";

when "001101101001101" => rgb <= "000000";

when "001101101001110" => rgb <= "100110";

when "001101101001111" => rgb <= "100110";

when "001101101010000" => rgb <= "100110";

when "001101101010001" => rgb <= "000000";

when "001101101010010" => rgb <= "000000";

when "001101101010101" => rgb <= "000000";

when "001101101010110" => rgb <= "000000";

when "001101101010111" => rgb <= "100110";

when "001101101011000" => rgb <= "100110";

when "001101101011001" => rgb <= "100110";

when "001101101011010" => rgb <= "000000";

when "001101101011101" => rgb <= "000000";

when "001101101011110" => rgb <= "100110";

when "001101101011111" => rgb <= "100110";

when "001101101100000" => rgb <= "100110";

when "001101101100001" => rgb <= "100110";

when "001101101100010" => rgb <= "100110";

when "001101101100011" => rgb <= "100110";

when "001101101100100" => rgb <= "100110";

when "001101101100101" => rgb <= "100110";

when "001101101100110" => rgb <= "000000";

when "001101101100111" => rgb <= "000000";

when "001110000110001" => rgb <= "000000";

when "001110000110010" => rgb <= "100110";

when "001110000110011" => rgb <= "100110";

when "001110000110100" => rgb <= "100110";

when "001110000110101" => rgb <= "100110";

when "001110000110110" => rgb <= "000000";

when "001110000111101" => rgb <= "000000";

when "001110000111110" => rgb <= "100110";

when "001110000111111" => rgb <= "100110";

when "001110001000000" => rgb <= "100110";

when "001110001000001" => rgb <= "000000";

when "001110001000010" => rgb <= "000000";

when "001110001000101" => rgb <= "000000";

when "001110001000110" => rgb <= "000000";

when "001110001000111" => rgb <= "100110";

when "001110001001000" => rgb <= "100110";

when "001110001001001" => rgb <= "100110";

when "001110001001010" => rgb <= "000000";

when "001110001001101" => rgb <= "000000";

when "001110001001110" => rgb <= "100110";

when "001110001001111" => rgb <= "100110";

when "001110001010000" => rgb <= "100110";

when "001110001010001" => rgb <= "100110";

when "001110001010010" => rgb <= "000000";

when "001110001010101" => rgb <= "000000";

when "001110001010110" => rgb <= "100110";

when "001110001010111" => rgb <= "100110";

when "001110001011000" => rgb <= "100110";

when "001110001011001" => rgb <= "100110";

when "001110001011010" => rgb <= "000000";

when "001110001011101" => rgb <= "000000";

when "001110001011110" => rgb <= "100110";

when "001110001011111" => rgb <= "100110";

when "001110001100000" => rgb <= "100110";

when "001110001100001" => rgb <= "000000";

when "001110001100010" => rgb <= "000000";

when "001110001100011" => rgb <= "100110";

when "001110001100100" => rgb <= "100110";

when "001110001100101" => rgb <= "100110";

when "001110001100110" => rgb <= "100110";

when "001110001100111" => rgb <= "000000";

when "001110001101000" => rgb <= "000000";

when "001110100110001" => rgb <= "000000";

when "001110100110010" => rgb <= "100110";

when "001110100110011" => rgb <= "100110";

when "001110100110100" => rgb <= "100110";

when "001110100110101" => rgb <= "100110";

when "001110100110110" => rgb <= "000000";

when "001110100111101" => rgb <= "000000";

when "001110100111110" => rgb <= "100110";

when "001110100111111" => rgb <= "100110";

when "001110101000000" => rgb <= "100110";

when "001110101000001" => rgb <= "100110";

when "001110101000010" => rgb <= "000000";

when "001110101000011" => rgb <= "000000";

when "001110101000100" => rgb <= "000000";

when "001110101000101" => rgb <= "000000";

when "001110101000110" => rgb <= "100110";

when "001110101000111" => rgb <= "100110";

when "001110101001000" => rgb <= "100110";

when "001110101001001" => rgb <= "100110";

when "001110101001010" => rgb <= "000000";

when "001110101001101" => rgb <= "000000";

when "001110101001110" => rgb <= "000000";

when "001110101001111" => rgb <= "100110";

when "001110101010000" => rgb <= "100110";

when "001110101010001" => rgb <= "100110";

when "001110101010010" => rgb <= "000000";

when "001110101010011" => rgb <= "000000";

when "001110101010100" => rgb <= "000000";

when "001110101010101" => rgb <= "000000";

when "001110101010110" => rgb <= "100110";

when "001110101010111" => rgb <= "100110";

when "001110101011000" => rgb <= "100110";

when "001110101011001" => rgb <= "000000";

when "001110101011010" => rgb <= "000000";

when "001110101011101" => rgb <= "000000";

when "001110101011110" => rgb <= "100110";

when "001110101011111" => rgb <= "100110";

when "001110101100000" => rgb <= "100110";

when "001110101100001" => rgb <= "000000";

when "001110101100011" => rgb <= "000000";

when "001110101100100" => rgb <= "100110";

when "001110101100101" => rgb <= "100110";

when "001110101100110" => rgb <= "100110";

when "001110101100111" => rgb <= "100110";

when "001110101101000" => rgb <= "000000";

when "001110101101001" => rgb <= "000000";

when "001111000110001" => rgb <= "000000";

when "001111000110010" => rgb <= "100110";

when "001111000110011" => rgb <= "100110";

when "001111000110100" => rgb <= "100110";

when "001111000110101" => rgb <= "100110";

when "001111000110110" => rgb <= "000000";

when "001111000111101" => rgb <= "000000";

when "001111000111110" => rgb <= "000000";

when "001111000111111" => rgb <= "100110";

when "001111001000000" => rgb <= "100110";

when "001111001000001" => rgb <= "100110";

when "001111001000010" => rgb <= "100110";

when "001111001000011" => rgb <= "100110";

when "001111001000100" => rgb <= "100110";

when "001111001000101" => rgb <= "100110";

when "001111001000110" => rgb <= "100110";

when "001111001000111" => rgb <= "100110";

when "001111001001000" => rgb <= "100110";

when "001111001001001" => rgb <= "000000";

when "001111001001010" => rgb <= "000000";

when "001111001001110" => rgb <= "000000";

when "001111001001111" => rgb <= "100110";

when "001111001010000" => rgb <= "100110";

when "001111001010001" => rgb <= "100110";

when "001111001010010" => rgb <= "100110";

when "001111001010011" => rgb <= "100110";

when "001111001010100" => rgb <= "100110";

when "001111001010101" => rgb <= "100110";

when "001111001010110" => rgb <= "100110";

when "001111001010111" => rgb <= "100110";

when "001111001011000" => rgb <= "100110";

when "001111001011001" => rgb <= "000000";

when "001111001011101" => rgb <= "000000";

when "001111001011110" => rgb <= "100110";

when "001111001011111" => rgb <= "100110";

when "001111001100000" => rgb <= "100110";

when "001111001100001" => rgb <= "000000";

when "001111001100011" => rgb <= "000000";

when "001111001100100" => rgb <= "000000";

when "001111001100101" => rgb <= "100110";

when "001111001100110" => rgb <= "100110";

when "001111001100111" => rgb <= "100110";

when "001111001101000" => rgb <= "100110";

when "001111001101001" => rgb <= "000000";

when "001111100110001" => rgb <= "000000";

when "001111100110010" => rgb <= "100110";

when "001111100110011" => rgb <= "100110";

when "001111100110100" => rgb <= "100110";

when "001111100110101" => rgb <= "100110";

when "001111100110110" => rgb <= "000000";

when "001111100111110" => rgb <= "000000";

when "001111100111111" => rgb <= "100110";

when "001111101000000" => rgb <= "100110";

when "001111101000001" => rgb <= "100110";

when "001111101000010" => rgb <= "100110";

when "001111101000011" => rgb <= "100110";

when "001111101000100" => rgb <= "100110";

when "001111101000101" => rgb <= "100110";

when "001111101000110" => rgb <= "100110";

when "001111101000111" => rgb <= "100110";

when "001111101001000" => rgb <= "100110";

when "001111101001001" => rgb <= "000000";

when "001111101001110" => rgb <= "000000";

when "001111101001111" => rgb <= "000000";

when "001111101010000" => rgb <= "100110";

when "001111101010001" => rgb <= "100110";

when "001111101010010" => rgb <= "100110";

when "001111101010011" => rgb <= "100110";

when "001111101010100" => rgb <= "100110";

when "001111101010101" => rgb <= "100110";

when "001111101010110" => rgb <= "100110";

when "001111101010111" => rgb <= "100110";

when "001111101011000" => rgb <= "000000";

when "001111101011001" => rgb <= "000000";

when "001111101011101" => rgb <= "000000";

when "001111101011110" => rgb <= "100110";

when "001111101011111" => rgb <= "100110";

when "001111101100000" => rgb <= "100110";

when "001111101100001" => rgb <= "000000";

when "001111101100100" => rgb <= "000000";

when "001111101100101" => rgb <= "000000";

when "001111101100110" => rgb <= "100110";

when "001111101100111" => rgb <= "100110";

when "001111101101000" => rgb <= "100110";

when "001111101101001" => rgb <= "000000";

when "010000000110001" => rgb <= "000000";

when "010000000110010" => rgb <= "100110";

when "010000000110011" => rgb <= "100110";

when "010000000110100" => rgb <= "100110";

when "010000000110101" => rgb <= "100110";

when "010000000110110" => rgb <= "000000";

when "010000000111110" => rgb <= "000000";

when "010000000111111" => rgb <= "000000";

when "010000001000000" => rgb <= "000000";

when "010000001000001" => rgb <= "100110";

when "010000001000010" => rgb <= "100110";

when "010000001000011" => rgb <= "100110";

when "010000001000100" => rgb <= "100110";

when "010000001000101" => rgb <= "100110";

when "010000001000110" => rgb <= "100110";

when "010000001000111" => rgb <= "000000";

when "010000001001000" => rgb <= "000000";

when "010000001001001" => rgb <= "000000";

when "010000001001111" => rgb <= "000000";

when "010000001010000" => rgb <= "100110";

when "010000001010001" => rgb <= "100110";

when "010000001010010" => rgb <= "100110";

when "010000001010011" => rgb <= "100110";

when "010000001010100" => rgb <= "100110";

when "010000001010101" => rgb <= "100110";

when "010000001010110" => rgb <= "100110";

when "010000001010111" => rgb <= "100110";

when "010000001011000" => rgb <= "000000";

when "010000001011101" => rgb <= "000000";

when "010000001011110" => rgb <= "100110";

when "010000001011111" => rgb <= "100110";

when "010000001100000" => rgb <= "100110";

when "010000001100001" => rgb <= "000000";

when "010000001100101" => rgb <= "000000";

when "010000001100110" => rgb <= "100110";

when "010000001100111" => rgb <= "100110";

when "010000001101000" => rgb <= "100110";

when "010000001101001" => rgb <= "000000";

when "010000100110001" => rgb <= "000000";

when "010000100110010" => rgb <= "000000";

when "010000100110011" => rgb <= "000000";

when "010000100110100" => rgb <= "000000";

when "010000100110101" => rgb <= "000000";

when "010000100110110" => rgb <= "000000";

when "010000101000000" => rgb <= "000000";

when "010000101000001" => rgb <= "000000";

when "010000101000010" => rgb <= "000000";

when "010000101000011" => rgb <= "000000";

when "010000101000100" => rgb <= "000000";

when "010000101000101" => rgb <= "000000";

when "010000101000110" => rgb <= "000000";

when "010000101000111" => rgb <= "000000";

when "010000101001111" => rgb <= "000000";

when "010000101010000" => rgb <= "000000";

when "010000101010001" => rgb <= "000000";

when "010000101010010" => rgb <= "000000";

when "010000101010011" => rgb <= "000000";

when "010000101010100" => rgb <= "000000";

when "010000101010101" => rgb <= "000000";

when "010000101010110" => rgb <= "000000";

when "010000101010111" => rgb <= "000000";

when "010000101011000" => rgb <= "000000";

when "010000101011101" => rgb <= "000000";

when "010000101011110" => rgb <= "000000";

when "010000101011111" => rgb <= "000000";

when "010000101100000" => rgb <= "000000";

when "010000101100001" => rgb <= "000000";

when "010000101100101" => rgb <= "000000";

when "010000101100110" => rgb <= "000000";

when "010000101100111" => rgb <= "000000";

when "010000101101000" => rgb <= "000000";

when "010000101101001" => rgb <= "000000";

when "010100000101110" => rgb <= "000000";

when "010100000101111" => rgb <= "000000";

when "010100000110000" => rgb <= "000000";

when "010100000110001" => rgb <= "000000";

when "010100000110010" => rgb <= "000000";

when "010100000110011" => rgb <= "000000";

when "010100000110100" => rgb <= "000000";

when "010100000110101" => rgb <= "000000";

when "010100000110110" => rgb <= "000000";

when "010100000110111" => rgb <= "000000";

when "010100000111000" => rgb <= "000000";

when "010100000111001" => rgb <= "000000";

when "010100000111010" => rgb <= "000000";

when "010100000111101" => rgb <= "000000";

when "010100000111110" => rgb <= "000000";

when "010100000111111" => rgb <= "000000";

when "010100001000000" => rgb <= "000000";

when "010100001000001" => rgb <= "000000";

when "010100001000110" => rgb <= "000000";

when "010100001000111" => rgb <= "000000";

when "010100001001000" => rgb <= "000000";

when "010100001001001" => rgb <= "000000";

when "010100001001010" => rgb <= "000000";

when "010100001001101" => rgb <= "000000";

when "010100001001110" => rgb <= "000000";

when "010100001001111" => rgb <= "000000";

when "010100001010000" => rgb <= "000000";

when "010100001010001" => rgb <= "000000";

when "010100001010010" => rgb <= "000000";

when "010100001010011" => rgb <= "000000";

when "010100001010100" => rgb <= "000000";

when "010100001010101" => rgb <= "000000";

when "010100001010110" => rgb <= "000000";

when "010100001010111" => rgb <= "000000";

when "010100001011100" => rgb <= "000000";

when "010100001011101" => rgb <= "000000";

when "010100001011110" => rgb <= "000000";

when "010100001011111" => rgb <= "000000";

when "010100001100000" => rgb <= "000000";

when "010100001100001" => rgb <= "000000";

when "010100001100100" => rgb <= "000000";

when "010100001100101" => rgb <= "000000";

when "010100001100110" => rgb <= "000000";

when "010100001100111" => rgb <= "000000";

when "010100001101000" => rgb <= "000000";

when "010100100101110" => rgb <= "000000";

when "010100100101111" => rgb <= "100110";

when "010100100110000" => rgb <= "100110";

when "010100100110001" => rgb <= "100110";

when "010100100110010" => rgb <= "100110";

when "010100100110011" => rgb <= "100110";

when "010100100110100" => rgb <= "100110";

when "010100100110101" => rgb <= "100110";

when "010100100110110" => rgb <= "100110";

when "010100100110111" => rgb <= "100110";

when "010100100111000" => rgb <= "100110";

when "010100100111001" => rgb <= "100110";

when "010100100111010" => rgb <= "000000";

when "010100100111101" => rgb <= "000000";

when "010100100111110" => rgb <= "100110";

when "010100100111111" => rgb <= "100110";

when "010100101000000" => rgb <= "100110";

when "010100101000001" => rgb <= "000000";

when "010100101000110" => rgb <= "000000";

when "010100101000111" => rgb <= "100110";

when "010100101001000" => rgb <= "100110";

when "010100101001001" => rgb <= "100110";

when "010100101001010" => rgb <= "000000";

when "010100101001101" => rgb <= "000000";

when "010100101001110" => rgb <= "100110";

when "010100101001111" => rgb <= "100110";

when "010100101010000" => rgb <= "100110";

when "010100101010001" => rgb <= "100110";

when "010100101010010" => rgb <= "100110";

when "010100101010011" => rgb <= "100110";

when "010100101010100" => rgb <= "100110";

when "010100101010101" => rgb <= "100110";

when "010100101010110" => rgb <= "100110";

when "010100101010111" => rgb <= "000000";

when "010100101011000" => rgb <= "000000";

when "010100101011001" => rgb <= "000000";

when "010100101011100" => rgb <= "000000";

when "010100101011101" => rgb <= "100110";

when "010100101011110" => rgb <= "100110";

when "010100101011111" => rgb <= "100110";

when "010100101100000" => rgb <= "100110";

when "010100101100001" => rgb <= "000000";

when "010100101100100" => rgb <= "000000";

when "010100101100101" => rgb <= "100110";

when "010100101100110" => rgb <= "100110";

when "010100101100111" => rgb <= "100110";

when "010100101101000" => rgb <= "000000";

when "010101000101110" => rgb <= "000000";

when "010101000101111" => rgb <= "100110";

when "010101000110000" => rgb <= "100110";

when "010101000110001" => rgb <= "100110";

when "010101000110010" => rgb <= "100110";

when "010101000110011" => rgb <= "100110";

when "010101000110100" => rgb <= "100110";

when "010101000110101" => rgb <= "100110";

when "010101000110110" => rgb <= "100110";

when "010101000110111" => rgb <= "100110";

when "010101000111000" => rgb <= "100110";

when "010101000111001" => rgb <= "100110";

when "010101000111010" => rgb <= "000000";

when "010101000111101" => rgb <= "000000";

when "010101000111110" => rgb <= "100110";

when "010101000111111" => rgb <= "100110";

when "010101001000000" => rgb <= "100110";

when "010101001000001" => rgb <= "000000";

when "010101001000110" => rgb <= "000000";

when "010101001000111" => rgb <= "100110";

when "010101001001000" => rgb <= "100110";

when "010101001001001" => rgb <= "100110";

when "010101001001010" => rgb <= "000000";

when "010101001001101" => rgb <= "000000";

when "010101001001110" => rgb <= "100110";

when "010101001001111" => rgb <= "100110";

when "010101001010000" => rgb <= "100110";

when "010101001010001" => rgb <= "100110";

when "010101001010010" => rgb <= "100110";

when "010101001010011" => rgb <= "100110";

when "010101001010100" => rgb <= "100110";

when "010101001010101" => rgb <= "100110";

when "010101001010110" => rgb <= "100110";

when "010101001010111" => rgb <= "100110";

when "010101001011000" => rgb <= "100110";

when "010101001011001" => rgb <= "000000";

when "010101001011100" => rgb <= "000000";

when "010101001011101" => rgb <= "100110";

when "010101001011110" => rgb <= "100110";

when "010101001011111" => rgb <= "100110";

when "010101001100000" => rgb <= "100110";

when "010101001100001" => rgb <= "000000";

when "010101001100010" => rgb <= "000000";

when "010101001100100" => rgb <= "000000";

when "010101001100101" => rgb <= "100110";

when "010101001100110" => rgb <= "100110";

when "010101001100111" => rgb <= "100110";

when "010101001101000" => rgb <= "000000";

when "010101100101110" => rgb <= "000000";

when "010101100101111" => rgb <= "100110";

when "010101100110000" => rgb <= "100110";

when "010101100110001" => rgb <= "100110";

when "010101100110010" => rgb <= "100110";

when "010101100110011" => rgb <= "100110";

when "010101100110100" => rgb <= "100110";

when "010101100110101" => rgb <= "100110";

when "010101100110110" => rgb <= "100110";

when "010101100110111" => rgb <= "100110";

when "010101100111000" => rgb <= "100110";

when "010101100111001" => rgb <= "100110";

when "010101100111010" => rgb <= "000000";

when "010101100111101" => rgb <= "000000";

when "010101100111110" => rgb <= "100110";

when "010101100111111" => rgb <= "100110";

when "010101101000000" => rgb <= "100110";

when "010101101000001" => rgb <= "000000";

when "010101101000110" => rgb <= "000000";

when "010101101000111" => rgb <= "100110";

when "010101101001000" => rgb <= "100110";

when "010101101001001" => rgb <= "100110";

when "010101101001010" => rgb <= "000000";

when "010101101001101" => rgb <= "000000";

when "010101101001110" => rgb <= "100110";

when "010101101001111" => rgb <= "100110";

when "010101101010000" => rgb <= "100110";

when "010101101010001" => rgb <= "000000";

when "010101101010010" => rgb <= "000000";

when "010101101010011" => rgb <= "000000";

when "010101101010100" => rgb <= "000000";

when "010101101010101" => rgb <= "000000";

when "010101101010110" => rgb <= "100110";

when "010101101010111" => rgb <= "100110";

when "010101101011000" => rgb <= "100110";

when "010101101011001" => rgb <= "000000";

when "010101101011100" => rgb <= "000000";

when "010101101011101" => rgb <= "100110";

when "010101101011110" => rgb <= "100110";

when "010101101011111" => rgb <= "100110";

when "010101101100000" => rgb <= "100110";

when "010101101100001" => rgb <= "100110";

when "010101101100010" => rgb <= "000000";

when "010101101100100" => rgb <= "000000";

when "010101101100101" => rgb <= "100110";

when "010101101100110" => rgb <= "100110";

when "010101101100111" => rgb <= "100110";

when "010101101101000" => rgb <= "000000";

when "010110000101110" => rgb <= "000000";

when "010110000101111" => rgb <= "000000";

when "010110000110000" => rgb <= "000000";

when "010110000110001" => rgb <= "000000";

when "010110000110010" => rgb <= "000000";

when "010110000110011" => rgb <= "100110";

when "010110000110100" => rgb <= "100110";

when "010110000110101" => rgb <= "100110";

when "010110000110110" => rgb <= "000000";

when "010110000110111" => rgb <= "000000";

when "010110000111000" => rgb <= "000000";

when "010110000111001" => rgb <= "000000";

when "010110000111010" => rgb <= "000000";

when "010110000111101" => rgb <= "000000";

when "010110000111110" => rgb <= "100110";

when "010110000111111" => rgb <= "100110";

when "010110001000000" => rgb <= "100110";

when "010110001000001" => rgb <= "000000";

when "010110001000110" => rgb <= "000000";

when "010110001000111" => rgb <= "100110";

when "010110001001000" => rgb <= "100110";

when "010110001001001" => rgb <= "100110";

when "010110001001010" => rgb <= "000000";

when "010110001001101" => rgb <= "000000";

when "010110001001110" => rgb <= "100110";

when "010110001001111" => rgb <= "100110";

when "010110001010000" => rgb <= "100110";

when "010110001010001" => rgb <= "000000";

when "010110001010101" => rgb <= "000000";

when "010110001010110" => rgb <= "100110";

when "010110001010111" => rgb <= "100110";

when "010110001011000" => rgb <= "100110";

when "010110001011001" => rgb <= "000000";

when "010110001011100" => rgb <= "000000";

when "010110001011101" => rgb <= "100110";

when "010110001011110" => rgb <= "100110";

when "010110001011111" => rgb <= "100110";

when "010110001100000" => rgb <= "100110";

when "010110001100001" => rgb <= "100110";

when "010110001100010" => rgb <= "000000";

when "010110001100011" => rgb <= "000000";

when "010110001100100" => rgb <= "000000";

when "010110001100101" => rgb <= "100110";

when "010110001100110" => rgb <= "100110";

when "010110001100111" => rgb <= "100110";

when "010110001101000" => rgb <= "000000";

when "010110100110010" => rgb <= "000000";

when "010110100110011" => rgb <= "100110";

when "010110100110100" => rgb <= "100110";

when "010110100110101" => rgb <= "100110";

when "010110100110110" => rgb <= "000000";

when "010110100111101" => rgb <= "000000";

when "010110100111110" => rgb <= "100110";

when "010110100111111" => rgb <= "100110";

when "010110101000000" => rgb <= "100110";

when "010110101000001" => rgb <= "000000";

when "010110101000110" => rgb <= "000000";

when "010110101000111" => rgb <= "100110";

when "010110101001000" => rgb <= "100110";

when "010110101001001" => rgb <= "100110";

when "010110101001010" => rgb <= "000000";

when "010110101001101" => rgb <= "000000";

when "010110101001110" => rgb <= "100110";

when "010110101001111" => rgb <= "100110";

when "010110101010000" => rgb <= "100110";

when "010110101010001" => rgb <= "000000";

when "010110101010101" => rgb <= "000000";

when "010110101010110" => rgb <= "100110";

when "010110101010111" => rgb <= "100110";

when "010110101011000" => rgb <= "100110";

when "010110101011001" => rgb <= "000000";

when "010110101011100" => rgb <= "000000";

when "010110101011101" => rgb <= "100110";

when "010110101011110" => rgb <= "100110";

when "010110101011111" => rgb <= "100110";

when "010110101100000" => rgb <= "100110";

when "010110101100001" => rgb <= "100110";

when "010110101100010" => rgb <= "100110";

when "010110101100011" => rgb <= "000000";

when "010110101100100" => rgb <= "000000";

when "010110101100101" => rgb <= "100110";

when "010110101100110" => rgb <= "100110";

when "010110101100111" => rgb <= "100110";

when "010110101101000" => rgb <= "000000";

when "010111000110010" => rgb <= "000000";

when "010111000110011" => rgb <= "100110";

when "010111000110100" => rgb <= "100110";

when "010111000110101" => rgb <= "100110";

when "010111000110110" => rgb <= "000000";

when "010111000111101" => rgb <= "000000";

when "010111000111110" => rgb <= "100110";

when "010111000111111" => rgb <= "100110";

when "010111001000000" => rgb <= "100110";

when "010111001000001" => rgb <= "000000";

when "010111001000110" => rgb <= "000000";

when "010111001000111" => rgb <= "100110";

when "010111001001000" => rgb <= "100110";

when "010111001001001" => rgb <= "100110";

when "010111001001010" => rgb <= "000000";

when "010111001001101" => rgb <= "000000";

when "010111001001110" => rgb <= "100110";

when "010111001001111" => rgb <= "100110";

when "010111001010000" => rgb <= "100110";

when "010111001010001" => rgb <= "000000";

when "010111001010100" => rgb <= "000000";

when "010111001010101" => rgb <= "000000";

when "010111001010110" => rgb <= "100110";

when "010111001010111" => rgb <= "100110";

when "010111001011000" => rgb <= "100110";

when "010111001011001" => rgb <= "000000";

when "010111001011100" => rgb <= "000000";

when "010111001011101" => rgb <= "100110";

when "010111001011110" => rgb <= "100110";

when "010111001011111" => rgb <= "100110";

when "010111001100000" => rgb <= "100110";

when "010111001100001" => rgb <= "100110";

when "010111001100010" => rgb <= "100110";

when "010111001100011" => rgb <= "100110";

when "010111001100100" => rgb <= "000000";

when "010111001100101" => rgb <= "100110";

when "010111001100110" => rgb <= "100110";

when "010111001100111" => rgb <= "100110";

when "010111001101000" => rgb <= "000000";

when "010111100110010" => rgb <= "000000";

when "010111100110011" => rgb <= "100110";

when "010111100110100" => rgb <= "100110";

when "010111100110101" => rgb <= "100110";

when "010111100110110" => rgb <= "000000";

when "010111100111101" => rgb <= "000000";

when "010111100111110" => rgb <= "100110";

when "010111100111111" => rgb <= "100110";

when "010111101000000" => rgb <= "100110";

when "010111101000001" => rgb <= "000000";

when "010111101000110" => rgb <= "000000";

when "010111101000111" => rgb <= "100110";

when "010111101001000" => rgb <= "100110";

when "010111101001001" => rgb <= "100110";

when "010111101001010" => rgb <= "000000";

when "010111101001101" => rgb <= "000000";

when "010111101001110" => rgb <= "100110";

when "010111101001111" => rgb <= "100110";

when "010111101010000" => rgb <= "100110";

when "010111101010001" => rgb <= "000000";

when "010111101010010" => rgb <= "000000";

when "010111101010011" => rgb <= "000000";

when "010111101010100" => rgb <= "000000";

when "010111101010101" => rgb <= "100110";

when "010111101010110" => rgb <= "100110";

when "010111101010111" => rgb <= "100110";

when "010111101011000" => rgb <= "100110";

when "010111101011001" => rgb <= "000000";

when "010111101011100" => rgb <= "000000";

when "010111101011101" => rgb <= "100110";

when "010111101011110" => rgb <= "100110";

when "010111101011111" => rgb <= "100110";

when "010111101100000" => rgb <= "100110";

when "010111101100001" => rgb <= "100110";

when "010111101100010" => rgb <= "100110";

when "010111101100011" => rgb <= "100110";

when "010111101100100" => rgb <= "100110";

when "010111101100101" => rgb <= "100110";

when "010111101100110" => rgb <= "100110";

when "010111101100111" => rgb <= "100110";

when "010111101101000" => rgb <= "000000";

when "011000000110010" => rgb <= "000000";

when "011000000110011" => rgb <= "100110";

when "011000000110100" => rgb <= "100110";

when "011000000110101" => rgb <= "100110";

when "011000000110110" => rgb <= "000000";

when "011000000111101" => rgb <= "000000";

when "011000000111110" => rgb <= "100110";

when "011000000111111" => rgb <= "100110";

when "011000001000000" => rgb <= "100110";

when "011000001000001" => rgb <= "000000";

when "011000001000110" => rgb <= "000000";

when "011000001000111" => rgb <= "100110";

when "011000001001000" => rgb <= "100110";

when "011000001001001" => rgb <= "100110";

when "011000001001010" => rgb <= "000000";

when "011000001001101" => rgb <= "000000";

when "011000001001110" => rgb <= "100110";

when "011000001001111" => rgb <= "100110";

when "011000001010000" => rgb <= "100110";

when "011000001010001" => rgb <= "100110";

when "011000001010010" => rgb <= "100110";

when "011000001010011" => rgb <= "100110";

when "011000001010100" => rgb <= "100110";

when "011000001010101" => rgb <= "100110";

when "011000001010110" => rgb <= "100110";

when "011000001010111" => rgb <= "000000";

when "011000001011000" => rgb <= "000000";

when "011000001011001" => rgb <= "000000";

when "011000001011100" => rgb <= "000000";

when "011000001011101" => rgb <= "100110";

when "011000001011110" => rgb <= "100110";

when "011000001011111" => rgb <= "100110";

when "011000001100000" => rgb <= "100110";

when "011000001100001" => rgb <= "100110";

when "011000001100010" => rgb <= "100110";

when "011000001100011" => rgb <= "100110";

when "011000001100100" => rgb <= "100110";

when "011000001100101" => rgb <= "100110";

when "011000001100110" => rgb <= "100110";

when "011000001100111" => rgb <= "100110";

when "011000001101000" => rgb <= "000000";

when "011000100110010" => rgb <= "000000";

when "011000100110011" => rgb <= "100110";

when "011000100110100" => rgb <= "100110";

when "011000100110101" => rgb <= "100110";

when "011000100110110" => rgb <= "000000";

when "011000100111101" => rgb <= "000000";

when "011000100111110" => rgb <= "100110";

when "011000100111111" => rgb <= "100110";

when "011000101000000" => rgb <= "100110";

when "011000101000001" => rgb <= "000000";

when "011000101000010" => rgb <= "000000";

when "011000101000101" => rgb <= "000000";

when "011000101000110" => rgb <= "000000";

when "011000101000111" => rgb <= "100110";

when "011000101001000" => rgb <= "100110";

when "011000101001001" => rgb <= "100110";

when "011000101001010" => rgb <= "000000";

when "011000101001101" => rgb <= "000000";

when "011000101001110" => rgb <= "100110";

when "011000101001111" => rgb <= "100110";

when "011000101010000" => rgb <= "100110";

when "011000101010001" => rgb <= "100110";

when "011000101010010" => rgb <= "100110";

when "011000101010011" => rgb <= "100110";

when "011000101010100" => rgb <= "100110";

when "011000101010101" => rgb <= "100110";

when "011000101010110" => rgb <= "000000";

when "011000101010111" => rgb <= "000000";

when "011000101011100" => rgb <= "000000";

when "011000101011101" => rgb <= "100110";

when "011000101011110" => rgb <= "100110";

when "011000101011111" => rgb <= "100110";

when "011000101100000" => rgb <= "000000";

when "011000101100001" => rgb <= "100110";

when "011000101100010" => rgb <= "100110";

when "011000101100011" => rgb <= "100110";

when "011000101100100" => rgb <= "100110";

when "011000101100101" => rgb <= "100110";

when "011000101100110" => rgb <= "100110";

when "011000101100111" => rgb <= "100110";

when "011000101101000" => rgb <= "000000";

when "011001000110010" => rgb <= "000000";

when "011001000110011" => rgb <= "100110";

when "011001000110100" => rgb <= "100110";

when "011001000110101" => rgb <= "100110";

when "011001000110110" => rgb <= "000000";

when "011001000111101" => rgb <= "000000";

when "011001000111110" => rgb <= "100110";

when "011001000111111" => rgb <= "100110";

when "011001001000000" => rgb <= "100110";

when "011001001000001" => rgb <= "100110";

when "011001001000010" => rgb <= "000000";

when "011001001000101" => rgb <= "000000";

when "011001001000110" => rgb <= "100110";

when "011001001000111" => rgb <= "100110";

when "011001001001000" => rgb <= "100110";

when "011001001001001" => rgb <= "100110";

when "011001001001010" => rgb <= "000000";

when "011001001001101" => rgb <= "000000";

when "011001001001110" => rgb <= "100110";

when "011001001001111" => rgb <= "100110";

when "011001001010000" => rgb <= "100110";

when "011001001010001" => rgb <= "000000";

when "011001001010010" => rgb <= "000000";

when "011001001010011" => rgb <= "100110";

when "011001001010100" => rgb <= "100110";

when "011001001010101" => rgb <= "100110";

when "011001001010110" => rgb <= "100110";

when "011001001010111" => rgb <= "000000";

when "011001001011000" => rgb <= "000000";

when "011001001011100" => rgb <= "000000";

when "011001001011101" => rgb <= "100110";

when "011001001011110" => rgb <= "100110";

when "011001001011111" => rgb <= "100110";

when "011001001100000" => rgb <= "000000";

when "011001001100001" => rgb <= "000000";

when "011001001100010" => rgb <= "100110";

when "011001001100011" => rgb <= "100110";

when "011001001100100" => rgb <= "100110";

when "011001001100101" => rgb <= "100110";

when "011001001100110" => rgb <= "100110";

when "011001001100111" => rgb <= "100110";

when "011001001101000" => rgb <= "000000";

when "011001100110010" => rgb <= "000000";

when "011001100110011" => rgb <= "100110";

when "011001100110100" => rgb <= "100110";

when "011001100110101" => rgb <= "100110";

when "011001100110110" => rgb <= "000000";

when "011001100111101" => rgb <= "000000";

when "011001100111110" => rgb <= "000000";

when "011001100111111" => rgb <= "100110";

when "011001101000000" => rgb <= "100110";

when "011001101000001" => rgb <= "100110";

when "011001101000010" => rgb <= "000000";

when "011001101000011" => rgb <= "000000";

when "011001101000100" => rgb <= "000000";

when "011001101000101" => rgb <= "000000";

when "011001101000110" => rgb <= "100110";

when "011001101000111" => rgb <= "100110";

when "011001101001000" => rgb <= "100110";

when "011001101001001" => rgb <= "000000";

when "011001101001010" => rgb <= "000000";

when "011001101001101" => rgb <= "000000";

when "011001101001110" => rgb <= "100110";

when "011001101001111" => rgb <= "100110";

when "011001101010000" => rgb <= "100110";

when "011001101010001" => rgb <= "000000";

when "011001101010011" => rgb <= "000000";

when "011001101010100" => rgb <= "100110";

when "011001101010101" => rgb <= "100110";

when "011001101010110" => rgb <= "100110";

when "011001101010111" => rgb <= "100110";

when "011001101011000" => rgb <= "000000";

when "011001101011001" => rgb <= "000000";

when "011001101011100" => rgb <= "000000";

when "011001101011101" => rgb <= "100110";

when "011001101011110" => rgb <= "100110";

when "011001101011111" => rgb <= "100110";

when "011001101100000" => rgb <= "000000";

when "011001101100001" => rgb <= "000000";

when "011001101100010" => rgb <= "000000";

when "011001101100011" => rgb <= "100110";

when "011001101100100" => rgb <= "100110";

when "011001101100101" => rgb <= "100110";

when "011001101100110" => rgb <= "100110";

when "011001101100111" => rgb <= "100110";

when "011001101101000" => rgb <= "000000";

when "011010000110010" => rgb <= "000000";

when "011010000110011" => rgb <= "100110";

when "011010000110100" => rgb <= "100110";

when "011010000110101" => rgb <= "100110";

when "011010000110110" => rgb <= "000000";

when "011010000111110" => rgb <= "000000";

when "011010000111111" => rgb <= "100110";

when "011010001000000" => rgb <= "100110";

when "011010001000001" => rgb <= "100110";

when "011010001000010" => rgb <= "100110";

when "011010001000011" => rgb <= "100110";

when "011010001000100" => rgb <= "100110";

when "011010001000101" => rgb <= "100110";

when "011010001000110" => rgb <= "100110";

when "011010001000111" => rgb <= "100110";

when "011010001001000" => rgb <= "100110";

when "011010001001001" => rgb <= "000000";

when "011010001001101" => rgb <= "000000";

when "011010001001110" => rgb <= "100110";

when "011010001001111" => rgb <= "100110";

when "011010001010000" => rgb <= "100110";

when "011010001010001" => rgb <= "000000";

when "011010001010011" => rgb <= "000000";

when "011010001010100" => rgb <= "000000";

when "011010001010101" => rgb <= "100110";

when "011010001010110" => rgb <= "100110";

when "011010001010111" => rgb <= "100110";

when "011010001011000" => rgb <= "100110";

when "011010001011001" => rgb <= "000000";

when "011010001011100" => rgb <= "000000";

when "011010001011101" => rgb <= "100110";

when "011010001011110" => rgb <= "100110";

when "011010001011111" => rgb <= "100110";

when "011010001100000" => rgb <= "000000";

when "011010001100010" => rgb <= "000000";

when "011010001100011" => rgb <= "100110";

when "011010001100100" => rgb <= "100110";

when "011010001100101" => rgb <= "100110";

when "011010001100110" => rgb <= "100110";

when "011010001100111" => rgb <= "100110";

when "011010001101000" => rgb <= "000000";

when "011010100110010" => rgb <= "000000";

when "011010100110011" => rgb <= "100110";

when "011010100110100" => rgb <= "100110";

when "011010100110101" => rgb <= "100110";

when "011010100110110" => rgb <= "000000";

when "011010100111110" => rgb <= "000000";

when "011010100111111" => rgb <= "000000";

when "011010101000000" => rgb <= "100110";

when "011010101000001" => rgb <= "100110";

when "011010101000010" => rgb <= "100110";

when "011010101000011" => rgb <= "100110";

when "011010101000100" => rgb <= "100110";

when "011010101000101" => rgb <= "100110";

when "011010101000110" => rgb <= "100110";

when "011010101000111" => rgb <= "100110";

when "011010101001000" => rgb <= "000000";

when "011010101001001" => rgb <= "000000";

when "011010101001101" => rgb <= "000000";

when "011010101001110" => rgb <= "100110";

when "011010101001111" => rgb <= "100110";

when "011010101010000" => rgb <= "100110";

when "011010101010001" => rgb <= "000000";

when "011010101010100" => rgb <= "000000";

when "011010101010101" => rgb <= "000000";

when "011010101010110" => rgb <= "100110";

when "011010101010111" => rgb <= "100110";

when "011010101011000" => rgb <= "100110";

when "011010101011001" => rgb <= "000000";

when "011010101011100" => rgb <= "000000";

when "011010101011101" => rgb <= "100110";

when "011010101011110" => rgb <= "100110";

when "011010101011111" => rgb <= "100110";

when "011010101100000" => rgb <= "000000";

when "011010101100010" => rgb <= "000000";

when "011010101100011" => rgb <= "000000";

when "011010101100100" => rgb <= "100110";

when "011010101100101" => rgb <= "100110";

when "011010101100110" => rgb <= "100110";

when "011010101100111" => rgb <= "100110";

when "011010101101000" => rgb <= "000000";

when "011011000110010" => rgb <= "000000";

when "011011000110011" => rgb <= "100110";

when "011011000110100" => rgb <= "100110";

when "011011000110101" => rgb <= "100110";

when "011011000110110" => rgb <= "000000";

when "011011000111111" => rgb <= "000000";

when "011011001000000" => rgb <= "100110";

when "011011001000001" => rgb <= "100110";

when "011011001000010" => rgb <= "100110";

when "011011001000011" => rgb <= "100110";

when "011011001000100" => rgb <= "100110";

when "011011001000101" => rgb <= "100110";

when "011011001000110" => rgb <= "100110";

when "011011001000111" => rgb <= "100110";

when "011011001001000" => rgb <= "000000";

when "011011001001101" => rgb <= "000000";

when "011011001001110" => rgb <= "100110";

when "011011001001111" => rgb <= "100110";

when "011011001010000" => rgb <= "100110";

when "011011001010001" => rgb <= "000000";

when "011011001010101" => rgb <= "000000";

when "011011001010110" => rgb <= "100110";

when "011011001010111" => rgb <= "100110";

when "011011001011000" => rgb <= "100110";

when "011011001011001" => rgb <= "000000";

when "011011001011100" => rgb <= "000000";

when "011011001011101" => rgb <= "100110";

when "011011001011110" => rgb <= "100110";

when "011011001011111" => rgb <= "100110";

when "011011001100000" => rgb <= "000000";

when "011011001100011" => rgb <= "000000";

when "011011001100100" => rgb <= "100110";

when "011011001100101" => rgb <= "100110";

when "011011001100110" => rgb <= "100110";

when "011011001100111" => rgb <= "100110";

when "011011001101000" => rgb <= "000000";

when "011011100110010" => rgb <= "000000";

when "011011100110011" => rgb <= "000000";

when "011011100110100" => rgb <= "000000";

when "011011100110101" => rgb <= "000000";

when "011011100110110" => rgb <= "000000";

when "011011100111111" => rgb <= "000000";

when "011011101000000" => rgb <= "000000";

when "011011101000001" => rgb <= "000000";

when "011011101000010" => rgb <= "000000";

when "011011101000011" => rgb <= "000000";

when "011011101000100" => rgb <= "000000";

when "011011101000101" => rgb <= "000000";

when "011011101000110" => rgb <= "000000";

when "011011101000111" => rgb <= "000000";

when "011011101001000" => rgb <= "000000";

when "011011101001101" => rgb <= "000000";

when "011011101001110" => rgb <= "000000";

when "011011101001111" => rgb <= "000000";

when "011011101010000" => rgb <= "000000";

when "011011101010001" => rgb <= "000000";

when "011011101010101" => rgb <= "000000";

when "011011101010110" => rgb <= "000000";

when "011011101010111" => rgb <= "000000";

when "011011101011000" => rgb <= "000000";

when "011011101011001" => rgb <= "000000";

when "011011101011100" => rgb <= "000000";

when "011011101011101" => rgb <= "000000";

when "011011101011110" => rgb <= "000000";

when "011011101011111" => rgb <= "000000";

when "011011101100000" => rgb <= "000000";

when "011011101100011" => rgb <= "000000";

when "011011101100100" => rgb <= "000000";

when "011011101100101" => rgb <= "000000";

when "011011101100110" => rgb <= "000000";

when "011011101100111" => rgb <= "000000";

when "011011101101000" => rgb <= "000000";
when others => rgb <= "111111"; --will update l8r
end case;
end if;
end process;
	addressOut <= address;
end;