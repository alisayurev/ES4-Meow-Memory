library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;


entity meow4 is --rom for the background
port(
    clk : in std_logic;
	address : in unsigned (14 downto 0); 
    rgb : out unsigned(5 downto 0)
);
end meow4;


architecture synth of meow4 is 

signal addressOut : unsigned(14 downto 0); 

begin
    process (clk) is begin
        if rising_edge(clk) then
            case addressOut is
                when "011010110000011" => rgb <= "000000";

when "011010110000100" => rgb <= "000000";

when "011010110000101" => rgb <= "000000";

when "011010110000110" => rgb <= "000000";

when "011010110000111" => rgb <= "000000";

when "011010110001000" => rgb <= "000000";

when "011010110001001" => rgb <= "000000";

when "011010110001010" => rgb <= "000000";

when "011010110001011" => rgb <= "000000";

when "011010110001100" => rgb <= "000000";

when "011010110001101" => rgb <= "000000";

when "011010110001110" => rgb <= "000000";

when "011010110001111" => rgb <= "000000";

when "011010110010000" => rgb <= "000000";

when "011010110010001" => rgb <= "000000";

when "011010110010010" => rgb <= "000000";

when "011010110010011" => rgb <= "000000";

when "011010110010100" => rgb <= "000000";

when "011010110010101" => rgb <= "000000";

when "011010110010110" => rgb <= "000000";

when "011010110010111" => rgb <= "000000";

when "011010110011000" => rgb <= "000000";

when "011010110011001" => rgb <= "000000";

when "011011010000010" => rgb <= "000000";

when "011011010000011" => rgb <= "111111";

when "011011010000100" => rgb <= "111111";

when "011011010000101" => rgb <= "111111";

when "011011010000110" => rgb <= "111111";

when "011011010000111" => rgb <= "111111";

when "011011010001000" => rgb <= "111111";

when "011011010001001" => rgb <= "111111";

when "011011010001010" => rgb <= "111111";

when "011011010001011" => rgb <= "111111";

when "011011010001100" => rgb <= "111111";

when "011011010001101" => rgb <= "111111";

when "011011010001110" => rgb <= "111111";

when "011011010001111" => rgb <= "111111";

when "011011010010000" => rgb <= "111111";

when "011011010010001" => rgb <= "111111";

when "011011010010010" => rgb <= "111111";

when "011011010010011" => rgb <= "111111";

when "011011010010100" => rgb <= "111111";

when "011011010010101" => rgb <= "111111";

when "011011010010110" => rgb <= "111111";

when "011011010010111" => rgb <= "111111";

when "011011010011000" => rgb <= "111111";

when "011011010011001" => rgb <= "111111";

when "011011010011010" => rgb <= "000000";

when "011011110000001" => rgb <= "000000";

when "011011110000010" => rgb <= "111111";

when "011011110000011" => rgb <= "111111";

when "011011110000100" => rgb <= "111111";

when "011011110000101" => rgb <= "111111";

when "011011110000110" => rgb <= "111111";

when "011011110000111" => rgb <= "111111";

when "011011110001000" => rgb <= "111111";

when "011011110001001" => rgb <= "111111";

when "011011110001010" => rgb <= "111111";

when "011011110001011" => rgb <= "111111";

when "011011110001100" => rgb <= "111111";

when "011011110001101" => rgb <= "111111";

when "011011110001110" => rgb <= "111111";

when "011011110001111" => rgb <= "111111";

when "011011110010000" => rgb <= "111111";

when "011011110010001" => rgb <= "111111";

when "011011110010010" => rgb <= "111111";

when "011011110010011" => rgb <= "111111";

when "011011110010100" => rgb <= "111111";

when "011011110010101" => rgb <= "111111";

when "011011110010110" => rgb <= "111111";

when "011011110010111" => rgb <= "111111";

when "011011110011000" => rgb <= "111111";

when "011011110011001" => rgb <= "111111";

when "011011110011010" => rgb <= "111111";

when "011011110011011" => rgb <= "000000";

when "011100010000001" => rgb <= "000000";

when "011100010000010" => rgb <= "111111";

when "011100010000011" => rgb <= "111111";

when "011100010000100" => rgb <= "111111";

when "011100010000101" => rgb <= "000000";

when "011100010000110" => rgb <= "000000";

when "011100010000111" => rgb <= "000000";

when "011100010001000" => rgb <= "000000";

when "011100010001001" => rgb <= "111111";

when "011100010001010" => rgb <= "111111";

when "011100010001011" => rgb <= "000000";

when "011100010001100" => rgb <= "000000";

when "011100010001101" => rgb <= "000000";

when "011100010001110" => rgb <= "111111";

when "011100010001111" => rgb <= "000000";

when "011100010010000" => rgb <= "000000";

when "011100010010001" => rgb <= "000000";

when "011100010010010" => rgb <= "111111";

when "011100010010011" => rgb <= "000000";

when "011100010010100" => rgb <= "111111";

when "011100010010101" => rgb <= "111111";

when "011100010010110" => rgb <= "111111";

when "011100010010111" => rgb <= "000000";

when "011100010011000" => rgb <= "111111";

when "011100010011001" => rgb <= "111111";

when "011100010011010" => rgb <= "111111";

when "011100010011011" => rgb <= "000000";

when "011100110000001" => rgb <= "000000";

when "011100110000010" => rgb <= "111111";

when "011100110000011" => rgb <= "111111";

when "011100110000100" => rgb <= "111111";

when "011100110000101" => rgb <= "000000";

when "011100110000110" => rgb <= "111111";

when "011100110000111" => rgb <= "000000";

when "011100110001000" => rgb <= "111111";

when "011100110001001" => rgb <= "000000";

when "011100110001010" => rgb <= "111111";

when "011100110001011" => rgb <= "000000";

when "011100110001100" => rgb <= "111111";

when "011100110001101" => rgb <= "111111";

when "011100110001110" => rgb <= "111111";

when "011100110001111" => rgb <= "000000";

when "011100110010000" => rgb <= "111111";

when "011100110010001" => rgb <= "000000";

when "011100110010010" => rgb <= "111111";

when "011100110010011" => rgb <= "000000";

when "011100110010100" => rgb <= "111111";

when "011100110010101" => rgb <= "111111";

when "011100110010110" => rgb <= "111111";

when "011100110010111" => rgb <= "000000";

when "011100110011000" => rgb <= "111111";

when "011100110011001" => rgb <= "111111";

when "011100110011010" => rgb <= "111111";

when "011100110011011" => rgb <= "000000";

when "011101010000001" => rgb <= "000000";

when "011101010000010" => rgb <= "111111";

when "011101010000011" => rgb <= "111111";

when "011101010000100" => rgb <= "111111";

when "011101010000101" => rgb <= "000000";

when "011101010000110" => rgb <= "111111";

when "011101010000111" => rgb <= "000000";

when "011101010001000" => rgb <= "111111";

when "011101010001001" => rgb <= "000000";

when "011101010001010" => rgb <= "111111";

when "011101010001011" => rgb <= "000000";

when "011101010001100" => rgb <= "000000";

when "011101010001101" => rgb <= "111111";

when "011101010001110" => rgb <= "111111";

when "011101010001111" => rgb <= "000000";

when "011101010010000" => rgb <= "111111";

when "011101010010001" => rgb <= "000000";

when "011101010010010" => rgb <= "111111";

when "011101010010011" => rgb <= "000000";

when "011101010010100" => rgb <= "111111";

when "011101010010101" => rgb <= "000000";

when "011101010010110" => rgb <= "111111";

when "011101010010111" => rgb <= "000000";

when "011101010011000" => rgb <= "111111";

when "011101010011001" => rgb <= "111111";

when "011101010011010" => rgb <= "111111";

when "011101010011011" => rgb <= "000000";

when "011101110000001" => rgb <= "000000";

when "011101110000010" => rgb <= "111111";

when "011101110000011" => rgb <= "111111";

when "011101110000100" => rgb <= "111111";

when "011101110000101" => rgb <= "000000";

when "011101110000110" => rgb <= "111111";

when "011101110000111" => rgb <= "000000";

when "011101110001000" => rgb <= "111111";

when "011101110001001" => rgb <= "000000";

when "011101110001010" => rgb <= "111111";

when "011101110001011" => rgb <= "000000";

when "011101110001100" => rgb <= "111111";

when "011101110001101" => rgb <= "111111";

when "011101110001110" => rgb <= "111111";

when "011101110001111" => rgb <= "000000";

when "011101110010000" => rgb <= "111111";

when "011101110010001" => rgb <= "000000";

when "011101110010010" => rgb <= "111111";

when "011101110010011" => rgb <= "000000";

when "011101110010100" => rgb <= "111111";

when "011101110010101" => rgb <= "000000";

when "011101110010110" => rgb <= "111111";

when "011101110010111" => rgb <= "000000";

when "011101110011000" => rgb <= "111111";

when "011101110011001" => rgb <= "111111";

when "011101110011010" => rgb <= "111111";

when "011101110011011" => rgb <= "000000";

when "011110010000001" => rgb <= "000000";

when "011110010000010" => rgb <= "111111";

when "011110010000011" => rgb <= "111111";

when "011110010000100" => rgb <= "111111";

when "011110010000101" => rgb <= "000000";

when "011110010000110" => rgb <= "111111";

when "011110010000111" => rgb <= "000000";

when "011110010001000" => rgb <= "111111";

when "011110010001001" => rgb <= "000000";

when "011110010001010" => rgb <= "111111";

when "011110010001011" => rgb <= "000000";

when "011110010001100" => rgb <= "000000";

when "011110010001101" => rgb <= "000000";

when "011110010001110" => rgb <= "111111";

when "011110010001111" => rgb <= "000000";

when "011110010010000" => rgb <= "000000";

when "011110010010001" => rgb <= "000000";

when "011110010010010" => rgb <= "111111";

when "011110010010011" => rgb <= "000000";

when "011110010010100" => rgb <= "000000";

when "011110010010101" => rgb <= "000000";

when "011110010010110" => rgb <= "000000";

when "011110010010111" => rgb <= "111111";

when "011110010011000" => rgb <= "111111";

when "011110010011001" => rgb <= "111111";

when "011110010011010" => rgb <= "111111";

when "011110010011011" => rgb <= "000000";

when "011110110000001" => rgb <= "000000";

when "011110110000010" => rgb <= "000000";

when "011110110000011" => rgb <= "111111";

when "011110110000100" => rgb <= "111111";

when "011110110000101" => rgb <= "111111";

when "011110110000110" => rgb <= "111111";

when "011110110000111" => rgb <= "111111";

when "011110110001000" => rgb <= "111111";

when "011110110001001" => rgb <= "111111";

when "011110110001010" => rgb <= "111111";

when "011110110001011" => rgb <= "111111";

when "011110110001100" => rgb <= "111111";

when "011110110001101" => rgb <= "111111";

when "011110110001110" => rgb <= "111111";

when "011110110001111" => rgb <= "111111";

when "011110110010000" => rgb <= "111111";

when "011110110010001" => rgb <= "111111";

when "011110110010010" => rgb <= "111111";

when "011110110010011" => rgb <= "111111";

when "011110110010100" => rgb <= "111111";

when "011110110010101" => rgb <= "111111";

when "011110110010110" => rgb <= "111111";

when "011110110010111" => rgb <= "111111";

when "011110110011000" => rgb <= "111111";

when "011110110011001" => rgb <= "111111";

when "011110110011010" => rgb <= "111111";

when "011110110011011" => rgb <= "000000";

when "011111010000010" => rgb <= "000000";

when "011111010000011" => rgb <= "111111";

when "011111010000100" => rgb <= "111111";

when "011111010000101" => rgb <= "111111";

when "011111010000110" => rgb <= "111111";

when "011111010000111" => rgb <= "111111";

when "011111010001000" => rgb <= "111111";

when "011111010001001" => rgb <= "111111";

when "011111010001010" => rgb <= "111111";

when "011111010001011" => rgb <= "111111";

when "011111010001100" => rgb <= "111111";

when "011111010001101" => rgb <= "111111";

when "011111010001110" => rgb <= "111111";

when "011111010001111" => rgb <= "111111";

when "011111010010000" => rgb <= "111111";

when "011111010010001" => rgb <= "111111";

when "011111010010010" => rgb <= "111111";

when "011111010010011" => rgb <= "111111";

when "011111010010100" => rgb <= "111111";

when "011111010010101" => rgb <= "111111";

when "011111010010110" => rgb <= "111111";

when "011111010010111" => rgb <= "111111";

when "011111010011000" => rgb <= "111111";

when "011111010011001" => rgb <= "111111";

when "011111010011010" => rgb <= "000000";

when "011111110000011" => rgb <= "000000";

when "011111110000100" => rgb <= "000000";

when "011111110000101" => rgb <= "000000";

when "011111110000110" => rgb <= "000000";

when "011111110000111" => rgb <= "111111";

when "011111110001000" => rgb <= "111111";

when "011111110001001" => rgb <= "111111";

when "011111110001010" => rgb <= "000000";

when "011111110001011" => rgb <= "000000";

when "011111110001100" => rgb <= "000000";

when "011111110001101" => rgb <= "000000";

when "011111110001110" => rgb <= "000000";

when "011111110001111" => rgb <= "000000";

when "011111110010000" => rgb <= "000000";

when "011111110010001" => rgb <= "000000";

when "011111110010010" => rgb <= "000000";

when "011111110010011" => rgb <= "000000";

when "011111110010100" => rgb <= "000000";

when "011111110010101" => rgb <= "000000";

when "011111110010110" => rgb <= "000000";

when "011111110010111" => rgb <= "000000";

when "011111110011000" => rgb <= "000000";

when "011111110011001" => rgb <= "000000";

when "100000010000110" => rgb <= "000000";

when "100000010000111" => rgb <= "111111";

when "100000010001000" => rgb <= "111111";

when "100000010001001" => rgb <= "111111";

when "100000010001010" => rgb <= "000000";

when "100000110000101" => rgb <= "000000";

when "100000110000110" => rgb <= "111111";

when "100000110000111" => rgb <= "111111";

when "100000110001000" => rgb <= "111111";

when "100000110001001" => rgb <= "000000";

when "100001010000101" => rgb <= "000000";

when "100001010000110" => rgb <= "111111";

when "100001010000111" => rgb <= "111111";

when "100001010001000" => rgb <= "000000";

when "100001110000101" => rgb <= "000000";

when "100001110000110" => rgb <= "000000";

when "100001110000111" => rgb <= "000000";
when others => rgb <= "110000"; --will update l8r
end case;
end if;
end process;
	addressOut <= address;
end;