library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;


entity pab is --rom for the background
port(
    clk : in std_logic;
	address : in unsigned (14 downto 0); 
    rgb : out unsigned(5 downto 0)
);
end pab;


architecture synth of pab is 

signal addressOut : unsigned(14 downto 0); 

begin
    process (clk) is begin
        if rising_edge(clk) then
            case addressOut is
                when "110011000011010" => rgb <= "000000";

when "110011000011011" => rgb <= "000000";

when "110011000011100" => rgb <= "000000";

when "110011000011110" => rgb <= "000000";

when "110011000011111" => rgb <= "000000";

when "110011000100010" => rgb <= "000000";

when "110011000100011" => rgb <= "000000";

when "110011000100100" => rgb <= "000000";

when "110011000100110" => rgb <= "000000";

when "110011000100111" => rgb <= "000000";

when "110011000101000" => rgb <= "000000";

when "110011000101010" => rgb <= "000000";

when "110011000101011" => rgb <= "000000";

when "110011000101100" => rgb <= "000000";

when "110011000110010" => rgb <= "000000";

when "110011000110011" => rgb <= "000000";

when "110011000110100" => rgb <= "000000";

when "110011000110110" => rgb <= "000000";

when "110011000111001" => rgb <= "000000";

when "110011000111011" => rgb <= "000000";

when "110011000111101" => rgb <= "000000";

when "110011001000011" => rgb <= "000000";

when "110011001000100" => rgb <= "000000";

when "110011001000111" => rgb <= "000000";

when "110011001001001" => rgb <= "000000";

when "110011001001011" => rgb <= "000000";

when "110011001001100" => rgb <= "000000";

when "110011001001101" => rgb <= "000000";

when "110011001001111" => rgb <= "000000";

when "110011001010000" => rgb <= "000000";

when "110011001010001" => rgb <= "000000";

when "110011001010011" => rgb <= "000000";

when "110011001010100" => rgb <= "000000";

when "110011001010101" => rgb <= "000000";

when "110011001010111" => rgb <= "000000";

when "110011001011010" => rgb <= "000000";

when "110011001100000" => rgb <= "000000";

when "110011001100001" => rgb <= "000000";

when "110011001100010" => rgb <= "000000";

when "110011001100100" => rgb <= "000000";

when "110011001100101" => rgb <= "000000";

when "110011001100110" => rgb <= "000000";

when "110011001101100" => rgb <= "000000";

when "110011001101101" => rgb <= "000000";

when "110011001110000" => rgb <= "000000";

when "110011001110001" => rgb <= "000000";

when "110011001110010" => rgb <= "000000";

when "110011001110100" => rgb <= "000000";

when "110011001110101" => rgb <= "000000";

when "110011001110110" => rgb <= "000000";

when "110011001111000" => rgb <= "000000";

when "110011001111010" => rgb <= "000000";

when "110011001111100" => rgb <= "000000";

when "110011001111101" => rgb <= "000000";

when "110011010000000" => rgb <= "000000";

when "110011010000011" => rgb <= "000000";

when "110011100011010" => rgb <= "000000";

when "110011100011100" => rgb <= "000000";

when "110011100011110" => rgb <= "000000";

when "110011100100000" => rgb <= "000000";

when "110011100100010" => rgb <= "000000";

when "110011100100110" => rgb <= "000000";

when "110011100101010" => rgb <= "000000";

when "110011100110010" => rgb <= "000000";

when "110011100110100" => rgb <= "000000";

when "110011100110110" => rgb <= "000000";

when "110011100110111" => rgb <= "000000";

when "110011100111001" => rgb <= "000000";

when "110011100111011" => rgb <= "000000";

when "110011100111101" => rgb <= "000000";

when "110011101000011" => rgb <= "000000";

when "110011101000101" => rgb <= "000000";

when "110011101000111" => rgb <= "000000";

when "110011101001001" => rgb <= "000000";

when "110011101001100" => rgb <= "000000";

when "110011101010000" => rgb <= "000000";

when "110011101010011" => rgb <= "000000";

when "110011101010101" => rgb <= "000000";

when "110011101010111" => rgb <= "000000";

when "110011101011000" => rgb <= "000000";

when "110011101011010" => rgb <= "000000";

when "110011101100001" => rgb <= "000000";

when "110011101100100" => rgb <= "000000";

when "110011101100110" => rgb <= "000000";

when "110011101101100" => rgb <= "000000";

when "110011101101110" => rgb <= "000000";

when "110011101110000" => rgb <= "000000";

when "110011101110101" => rgb <= "000000";

when "110011101111000" => rgb <= "000000";

when "110011101111010" => rgb <= "000000";

when "110011101111100" => rgb <= "000000";

when "110011101111110" => rgb <= "000000";

when "110011110000000" => rgb <= "000000";

when "110011110000001" => rgb <= "000000";

when "110011110000011" => rgb <= "000000";

when "110100000011010" => rgb <= "000000";

when "110100000011011" => rgb <= "000000";

when "110100000011100" => rgb <= "000000";

when "110100000011110" => rgb <= "000000";

when "110100000100000" => rgb <= "000000";

when "110100000100010" => rgb <= "000000";

when "110100000100011" => rgb <= "000000";

when "110100000100110" => rgb <= "000000";

when "110100000100111" => rgb <= "000000";

when "110100000101000" => rgb <= "000000";

when "110100000101010" => rgb <= "000000";

when "110100000101011" => rgb <= "000000";

when "110100000101100" => rgb <= "000000";

when "110100000110010" => rgb <= "000000";

when "110100000110011" => rgb <= "000000";

when "110100000110100" => rgb <= "000000";

when "110100000110110" => rgb <= "000000";

when "110100000111000" => rgb <= "000000";

when "110100000111001" => rgb <= "000000";

when "110100000111011" => rgb <= "000000";

when "110100000111101" => rgb <= "000000";

when "110100001000011" => rgb <= "000000";

when "110100001000100" => rgb <= "000000";

when "110100001000111" => rgb <= "000000";

when "110100001001001" => rgb <= "000000";

when "110100001001100" => rgb <= "000000";

when "110100001010000" => rgb <= "000000";

when "110100001010011" => rgb <= "000000";

when "110100001010101" => rgb <= "000000";

when "110100001010111" => rgb <= "000000";

when "110100001011001" => rgb <= "000000";

when "110100001011010" => rgb <= "000000";

when "110100001100001" => rgb <= "000000";

when "110100001100100" => rgb <= "000000";

when "110100001100110" => rgb <= "000000";

when "110100001101100" => rgb <= "000000";

when "110100001101110" => rgb <= "000000";

when "110100001110000" => rgb <= "000000";

when "110100001110001" => rgb <= "000000";

when "110100001110101" => rgb <= "000000";

when "110100001111000" => rgb <= "000000";

when "110100001111010" => rgb <= "000000";

when "110100001111100" => rgb <= "000000";

when "110100001111110" => rgb <= "000000";

when "110100010000000" => rgb <= "000000";

when "110100010000010" => rgb <= "000000";

when "110100010000011" => rgb <= "000000";

when "110100100011010" => rgb <= "000000";

when "110100100011110" => rgb <= "000000";

when "110100100011111" => rgb <= "000000";

when "110100100100010" => rgb <= "000000";

when "110100100101000" => rgb <= "000000";

when "110100100101100" => rgb <= "000000";

when "110100100110010" => rgb <= "000000";

when "110100100110100" => rgb <= "000000";

when "110100100110110" => rgb <= "000000";

when "110100100111001" => rgb <= "000000";

when "110100100111100" => rgb <= "000000";

when "110100101000011" => rgb <= "000000";

when "110100101000101" => rgb <= "000000";

when "110100101000111" => rgb <= "000000";

when "110100101001001" => rgb <= "000000";

when "110100101001100" => rgb <= "000000";

when "110100101010000" => rgb <= "000000";

when "110100101010011" => rgb <= "000000";

when "110100101010101" => rgb <= "000000";

when "110100101010111" => rgb <= "000000";

when "110100101011010" => rgb <= "000000";

when "110100101100001" => rgb <= "000000";

when "110100101100100" => rgb <= "000000";

when "110100101100110" => rgb <= "000000";

when "110100101101100" => rgb <= "000000";

when "110100101101101" => rgb <= "000000";

when "110100101110000" => rgb <= "000000";

when "110100101110101" => rgb <= "000000";

when "110100101111000" => rgb <= "000000";

when "110100101111010" => rgb <= "000000";

when "110100101111100" => rgb <= "000000";

when "110100101111101" => rgb <= "000000";

when "110100110000000" => rgb <= "000000";

when "110100110000011" => rgb <= "000000";

when "110101000011010" => rgb <= "000000";

when "110101000011110" => rgb <= "000000";

when "110101000100000" => rgb <= "000000";

when "110101000100010" => rgb <= "000000";

when "110101000100011" => rgb <= "000000";

when "110101000100100" => rgb <= "000000";

when "110101000100110" => rgb <= "000000";

when "110101000100111" => rgb <= "000000";

when "110101000101000" => rgb <= "000000";

when "110101000101010" => rgb <= "000000";

when "110101000101011" => rgb <= "000000";

when "110101000101100" => rgb <= "000000";

when "110101000110010" => rgb <= "000000";

when "110101000110100" => rgb <= "000000";

when "110101000110110" => rgb <= "000000";

when "110101000111001" => rgb <= "000000";

when "110101000111100" => rgb <= "000000";

when "110101001000011" => rgb <= "000000";

when "110101001000100" => rgb <= "000000";

when "110101001000101" => rgb <= "000000";

when "110101001000111" => rgb <= "000000";

when "110101001001000" => rgb <= "000000";

when "110101001001001" => rgb <= "000000";

when "110101001001100" => rgb <= "000000";

when "110101001010000" => rgb <= "000000";

when "110101001010011" => rgb <= "000000";

when "110101001010100" => rgb <= "000000";

when "110101001010101" => rgb <= "000000";

when "110101001010111" => rgb <= "000000";

when "110101001011010" => rgb <= "000000";

when "110101001100001" => rgb <= "000000";

when "110101001100100" => rgb <= "000000";

when "110101001100101" => rgb <= "000000";

when "110101001100110" => rgb <= "000000";

when "110101001101100" => rgb <= "000000";

when "110101001101110" => rgb <= "000000";

when "110101001110000" => rgb <= "000000";

when "110101001110001" => rgb <= "000000";

when "110101001110010" => rgb <= "000000";

when "110101001110101" => rgb <= "000000";

when "110101001111000" => rgb <= "000000";

when "110101001111001" => rgb <= "000000";

when "110101001111010" => rgb <= "000000";

when "110101001111100" => rgb <= "000000";

when "110101001111110" => rgb <= "000000";

when "110101010000000" => rgb <= "000000";

when "110101010000011" => rgb <= "000000";
when others => rgb <= "111111"; --will update l8r
end case;
end if;
end process;
	addressOut <= address;
end;