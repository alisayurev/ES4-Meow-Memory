library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;


entity meow2 is --rom for the background
port(
    clk : in std_logic;
	address : in unsigned (14 downto 0); 
    rgb : out unsigned(5 downto 0)
);
end meow2;


architecture synth of meow2 is 

signal addressOut : unsigned(14 downto 0); 

begin
    process (clk) is begin
        if rising_edge(clk) then
            case addressOut is
                when "011010100110111" => rgb <= "000000";

                when "011010100111000" => rgb <= "000000";
                
                when "011010100111001" => rgb <= "000000";
                
                when "011010100111010" => rgb <= "000000";
                
                when "011010100111011" => rgb <= "000000";
                
                when "011010100111100" => rgb <= "000000";
                
                when "011010100111101" => rgb <= "000000";
                
                when "011010100111110" => rgb <= "000000";
                
                when "011010100111111" => rgb <= "000000";
                
                when "011010101000000" => rgb <= "000000";
                
                when "011010101000001" => rgb <= "000000";
                
                when "011010101000010" => rgb <= "000000";
                
                when "011010101000011" => rgb <= "000000";
                
                when "011010101000100" => rgb <= "000000";
                
                when "011010101000101" => rgb <= "000000";
                
                when "011010101000110" => rgb <= "000000";
                
                when "011010101000111" => rgb <= "000000";
                
                when "011010101001000" => rgb <= "000000";
                
                when "011010101001001" => rgb <= "000000";
                
                when "011010101001010" => rgb <= "000000";
                
                when "011010101001011" => rgb <= "000000";
                
                when "011010101001100" => rgb <= "000000";
                
                when "011010101001101" => rgb <= "000000";
                
                when "011011000110110" => rgb <= "000000";
                
                when "011011000110111" => rgb <= "111111";
                
                when "011011000111000" => rgb <= "111111";
                
                when "011011000111001" => rgb <= "111111";
                
                when "011011000111010" => rgb <= "111111";
                
                when "011011000111011" => rgb <= "111111";
                
                when "011011000111100" => rgb <= "111111";
                
                when "011011000111101" => rgb <= "111111";
                
                when "011011000111110" => rgb <= "111111";
                
                when "011011000111111" => rgb <= "111111";
                
                when "011011001000000" => rgb <= "111111";
                
                when "011011001000001" => rgb <= "111111";
                
                when "011011001000010" => rgb <= "111111";
                
                when "011011001000011" => rgb <= "111111";
                
                when "011011001000100" => rgb <= "111111";
                
                when "011011001000101" => rgb <= "111111";
                
                when "011011001000110" => rgb <= "111111";
                
                when "011011001000111" => rgb <= "111111";
                
                when "011011001001000" => rgb <= "111111";
                
                when "011011001001001" => rgb <= "111111";
                
                when "011011001001010" => rgb <= "111111";
                
                when "011011001001011" => rgb <= "111111";
                
                when "011011001001100" => rgb <= "111111";
                
                when "011011001001101" => rgb <= "111111";
                
                when "011011001001110" => rgb <= "000000";
                
                when "011011100110101" => rgb <= "000000";
                
                when "011011100110110" => rgb <= "111111";
                
                when "011011100110111" => rgb <= "111111";
                
                when "011011100111000" => rgb <= "111111";
                
                when "011011100111001" => rgb <= "111111";
                
                when "011011100111010" => rgb <= "111111";
                
                when "011011100111011" => rgb <= "111111";
                
                when "011011100111100" => rgb <= "111111";
                
                when "011011100111101" => rgb <= "111111";
                
                when "011011100111110" => rgb <= "111111";
                
                when "011011100111111" => rgb <= "111111";
                
                when "011011101000000" => rgb <= "111111";
                
                when "011011101000001" => rgb <= "111111";
                
                when "011011101000010" => rgb <= "111111";
                
                when "011011101000011" => rgb <= "111111";
                
                when "011011101000100" => rgb <= "111111";
                
                when "011011101000101" => rgb <= "111111";
                
                when "011011101000110" => rgb <= "111111";
                
                when "011011101000111" => rgb <= "111111";
                
                when "011011101001000" => rgb <= "111111";
                
                when "011011101001001" => rgb <= "111111";
                
                when "011011101001010" => rgb <= "111111";
                
                when "011011101001011" => rgb <= "111111";
                
                when "011011101001100" => rgb <= "111111";
                
                when "011011101001101" => rgb <= "111111";
                
                when "011011101001110" => rgb <= "111111";
                
                when "011011101001111" => rgb <= "000000";
                
                when "011100000110101" => rgb <= "000000";
                
                when "011100000110110" => rgb <= "111111";
                
                when "011100000110111" => rgb <= "111111";
                
                when "011100000111000" => rgb <= "111111";
                
                when "011100000111001" => rgb <= "000000";
                
                when "011100000111010" => rgb <= "000000";
                
                when "011100000111011" => rgb <= "000000";
                
                when "011100000111100" => rgb <= "000000";
                
                when "011100000111101" => rgb <= "111111";
                
                when "011100000111110" => rgb <= "111111";
                
                when "011100000111111" => rgb <= "000000";
                
                when "011100001000000" => rgb <= "000000";
                
                when "011100001000001" => rgb <= "000000";
                
                when "011100001000010" => rgb <= "111111";
                
                when "011100001000011" => rgb <= "000000";
                
                when "011100001000100" => rgb <= "000000";
                
                when "011100001000101" => rgb <= "000000";
                
                when "011100001000110" => rgb <= "111111";
                
                when "011100001000111" => rgb <= "000000";
                
                when "011100001001000" => rgb <= "111111";
                
                when "011100001001001" => rgb <= "111111";
                
                when "011100001001010" => rgb <= "111111";
                
                when "011100001001011" => rgb <= "000000";
                
                when "011100001001100" => rgb <= "111111";
                
                when "011100001001101" => rgb <= "111111";
                
                when "011100001001110" => rgb <= "111111";
                
                when "011100001001111" => rgb <= "000000";
                
                when "011100100110101" => rgb <= "000000";
                
                when "011100100110110" => rgb <= "111111";
                
                when "011100100110111" => rgb <= "111111";
                
                when "011100100111000" => rgb <= "111111";
                
                when "011100100111001" => rgb <= "000000";
                
                when "011100100111010" => rgb <= "111111";
                
                when "011100100111011" => rgb <= "000000";
                
                when "011100100111100" => rgb <= "111111";
                
                when "011100100111101" => rgb <= "000000";
                
                when "011100100111110" => rgb <= "111111";
                
                when "011100100111111" => rgb <= "000000";
                
                when "011100101000000" => rgb <= "111111";
                
                when "011100101000001" => rgb <= "111111";
                
                when "011100101000010" => rgb <= "111111";
                
                when "011100101000011" => rgb <= "000000";
                
                when "011100101000100" => rgb <= "111111";
                
                when "011100101000101" => rgb <= "000000";
                
                when "011100101000110" => rgb <= "111111";
                
                when "011100101000111" => rgb <= "000000";
                
                when "011100101001000" => rgb <= "111111";
                
                when "011100101001001" => rgb <= "111111";
                
                when "011100101001010" => rgb <= "111111";
                
                when "011100101001011" => rgb <= "000000";
                
                when "011100101001100" => rgb <= "111111";
                
                when "011100101001101" => rgb <= "111111";
                
                when "011100101001110" => rgb <= "111111";
                
                when "011100101001111" => rgb <= "000000";
                
                when "011101000110101" => rgb <= "000000";
                
                when "011101000110110" => rgb <= "111111";
                
                when "011101000110111" => rgb <= "111111";
                
                when "011101000111000" => rgb <= "111111";
                
                when "011101000111001" => rgb <= "000000";
                
                when "011101000111010" => rgb <= "111111";
                
                when "011101000111011" => rgb <= "000000";
                
                when "011101000111100" => rgb <= "111111";
                
                when "011101000111101" => rgb <= "000000";
                
                when "011101000111110" => rgb <= "111111";
                
                when "011101000111111" => rgb <= "000000";
                
                when "011101001000000" => rgb <= "000000";
                
                when "011101001000001" => rgb <= "111111";
                
                when "011101001000010" => rgb <= "111111";
                
                when "011101001000011" => rgb <= "000000";
                
                when "011101001000100" => rgb <= "111111";
                
                when "011101001000101" => rgb <= "000000";
                
                when "011101001000110" => rgb <= "111111";
                
                when "011101001000111" => rgb <= "000000";
                
                when "011101001001000" => rgb <= "111111";
                
                when "011101001001001" => rgb <= "000000";
                
                when "011101001001010" => rgb <= "111111";
                
                when "011101001001011" => rgb <= "000000";
                
                when "011101001001100" => rgb <= "111111";
                
                when "011101001001101" => rgb <= "111111";
                
                when "011101001001110" => rgb <= "111111";
                
                when "011101001001111" => rgb <= "000000";
                
                when "011101100110101" => rgb <= "000000";
                
                when "011101100110110" => rgb <= "111111";
                
                when "011101100110111" => rgb <= "111111";
                
                when "011101100111000" => rgb <= "111111";
                
                when "011101100111001" => rgb <= "000000";
                
                when "011101100111010" => rgb <= "111111";
                
                when "011101100111011" => rgb <= "000000";
                
                when "011101100111100" => rgb <= "111111";
                
                when "011101100111101" => rgb <= "000000";
                
                when "011101100111110" => rgb <= "111111";
                
                when "011101100111111" => rgb <= "000000";
                
                when "011101101000000" => rgb <= "111111";
                
                when "011101101000001" => rgb <= "111111";
                
                when "011101101000010" => rgb <= "111111";
                
                when "011101101000011" => rgb <= "000000";
                
                when "011101101000100" => rgb <= "111111";
                
                when "011101101000101" => rgb <= "000000";
                
                when "011101101000110" => rgb <= "111111";
                
                when "011101101000111" => rgb <= "000000";
                
                when "011101101001000" => rgb <= "111111";
                
                when "011101101001001" => rgb <= "000000";
                
                when "011101101001010" => rgb <= "111111";
                
                when "011101101001011" => rgb <= "000000";
                
                when "011101101001100" => rgb <= "111111";
                
                when "011101101001101" => rgb <= "111111";
                
                when "011101101001110" => rgb <= "111111";
                
                when "011101101001111" => rgb <= "000000";
                
                when "011110000110101" => rgb <= "000000";
                
                when "011110000110110" => rgb <= "111111";
                
                when "011110000110111" => rgb <= "111111";
                
                when "011110000111000" => rgb <= "111111";
                
                when "011110000111001" => rgb <= "000000";
                
                when "011110000111010" => rgb <= "111111";
                
                when "011110000111011" => rgb <= "000000";
                
                when "011110000111100" => rgb <= "111111";
                
                when "011110000111101" => rgb <= "000000";
                
                when "011110000111110" => rgb <= "111111";
                
                when "011110000111111" => rgb <= "000000";
                
                when "011110001000000" => rgb <= "000000";
                
                when "011110001000001" => rgb <= "000000";
                
                when "011110001000010" => rgb <= "111111";
                
                when "011110001000011" => rgb <= "000000";
                
                when "011110001000100" => rgb <= "000000";
                
                when "011110001000101" => rgb <= "000000";
                
                when "011110001000110" => rgb <= "111111";
                
                when "011110001000111" => rgb <= "000000";
                
                when "011110001001000" => rgb <= "000000";
                
                when "011110001001001" => rgb <= "000000";
                
                when "011110001001010" => rgb <= "000000";
                
                when "011110001001011" => rgb <= "111111";
                
                when "011110001001100" => rgb <= "111111";
                
                when "011110001001101" => rgb <= "111111";
                
                when "011110001001110" => rgb <= "111111";
                
                when "011110001001111" => rgb <= "000000";
                
                when "011110100110101" => rgb <= "000000";
                
                when "011110100110110" => rgb <= "000000";
                
                when "011110100110111" => rgb <= "111111";
                
                when "011110100111000" => rgb <= "111111";
                
                when "011110100111001" => rgb <= "111111";
                
                when "011110100111010" => rgb <= "111111";
                
                when "011110100111011" => rgb <= "111111";
                
                when "011110100111100" => rgb <= "111111";
                
                when "011110100111101" => rgb <= "111111";
                
                when "011110100111110" => rgb <= "111111";
                
                when "011110100111111" => rgb <= "111111";
                
                when "011110101000000" => rgb <= "111111";
                
                when "011110101000001" => rgb <= "111111";
                
                when "011110101000010" => rgb <= "111111";
                
                when "011110101000011" => rgb <= "111111";
                
                when "011110101000100" => rgb <= "111111";
                
                when "011110101000101" => rgb <= "111111";
                
                when "011110101000110" => rgb <= "111111";
                
                when "011110101000111" => rgb <= "111111";
                
                when "011110101001000" => rgb <= "111111";
                
                when "011110101001001" => rgb <= "111111";
                
                when "011110101001010" => rgb <= "111111";
                
                when "011110101001011" => rgb <= "111111";
                
                when "011110101001100" => rgb <= "111111";
                
                when "011110101001101" => rgb <= "111111";
                
                when "011110101001110" => rgb <= "111111";
                
                when "011110101001111" => rgb <= "000000";
                
                when "011111000110110" => rgb <= "000000";
                
                when "011111000110111" => rgb <= "111111";
                
                when "011111000111000" => rgb <= "111111";
                
                when "011111000111001" => rgb <= "111111";
                
                when "011111000111010" => rgb <= "111111";
                
                when "011111000111011" => rgb <= "111111";
                
                when "011111000111100" => rgb <= "111111";
                
                when "011111000111101" => rgb <= "111111";
                
                when "011111000111110" => rgb <= "111111";
                
                when "011111000111111" => rgb <= "111111";
                
                when "011111001000000" => rgb <= "111111";
                
                when "011111001000001" => rgb <= "111111";
                
                when "011111001000010" => rgb <= "111111";
                
                when "011111001000011" => rgb <= "111111";
                
                when "011111001000100" => rgb <= "111111";
                
                when "011111001000101" => rgb <= "111111";
                
                when "011111001000110" => rgb <= "111111";
                
                when "011111001000111" => rgb <= "111111";
                
                when "011111001001000" => rgb <= "111111";
                
                when "011111001001001" => rgb <= "111111";
                
                when "011111001001010" => rgb <= "111111";
                
                when "011111001001011" => rgb <= "111111";
                
                when "011111001001100" => rgb <= "111111";
                
                when "011111001001101" => rgb <= "111111";
                
                when "011111001001110" => rgb <= "000000";
                
                when "011111100110111" => rgb <= "000000";
                
                when "011111100111000" => rgb <= "000000";
                
                when "011111100111001" => rgb <= "000000";
                
                when "011111100111010" => rgb <= "000000";
                
                when "011111100111011" => rgb <= "111111";
                
                when "011111100111100" => rgb <= "111111";
                
                when "011111100111101" => rgb <= "111111";
                
                when "011111100111110" => rgb <= "000000";
                
                when "011111100111111" => rgb <= "000000";
                
                when "011111101000000" => rgb <= "000000";
                
                when "011111101000001" => rgb <= "000000";
                
                when "011111101000010" => rgb <= "000000";
                
                when "011111101000011" => rgb <= "000000";
                
                when "011111101000100" => rgb <= "000000";
                
                when "011111101000101" => rgb <= "000000";
                
                when "011111101000110" => rgb <= "000000";
                
                when "011111101000111" => rgb <= "000000";
                
                when "011111101001000" => rgb <= "000000";
                
                when "011111101001001" => rgb <= "000000";
                
                when "011111101001010" => rgb <= "000000";
                
                when "011111101001011" => rgb <= "000000";
                
                when "011111101001100" => rgb <= "000000";
                
                when "011111101001101" => rgb <= "000000";
                
                when "100000000111010" => rgb <= "000000";
                
                when "100000000111011" => rgb <= "111111";
                
                when "100000000111100" => rgb <= "111111";
                
                when "100000000111101" => rgb <= "111111";
                
                when "100000000111110" => rgb <= "000000";
                
                when "100000100111001" => rgb <= "000000";
                
                when "100000100111010" => rgb <= "111111";
                
                when "100000100111011" => rgb <= "111111";
                
                when "100000100111100" => rgb <= "111111";
                
                when "100000100111101" => rgb <= "000000";
                
                when "100001000111001" => rgb <= "000000";
                
                when "100001000111010" => rgb <= "111111";
                
                when "100001000111011" => rgb <= "111111";
                
                when "100001000111100" => rgb <= "000000";
                
                when "100001100111001" => rgb <= "000000";
                
                when "100001100111010" => rgb <= "000000";
                
                when "100001100111011" => rgb <= "000000";
                when others => rgb <= "110000"; --will update l8r
end case;
end if;
end process;
	addressOut <= address;
end; 