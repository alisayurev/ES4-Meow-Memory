library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;


entity gameover is 
port(
    clk : in std_logic;
	address : in unsigned (14 downto 0); 
    rgb : out unsigned(5 downto 0)
);
end gameover;


architecture synth of gameover is 

signal addressOut : unsigned(14 downto 0); 

begin
    process (clk) is begin
        if rising_edge(clk) then
            case addressOut is
		when "000111000010101" => rgb <= "000000";
		when "000111000010110" => rgb <= "000000";
		when "000111000010111" => rgb <= "000000";
		when "000111000011000" => rgb <= "000000";
		when "000111000011001" => rgb <= "000000";
		when "000111000011010" => rgb <= "000000";
		when "000111000011011" => rgb <= "000000";
		when "000111000011100" => rgb <= "000000";
		when "000111000011101" => rgb <= "000000";
		when "000111000011110" => rgb <= "000000";
		when "000111000100011" => rgb <= "000000";
		when "000111000100100" => rgb <= "000000";
		when "000111000100101" => rgb <= "000000";
		when "000111000100110" => rgb <= "000000";
		when "000111000100111" => rgb <= "000000";
		when "000111000101000" => rgb <= "000000";
		when "000111000101001" => rgb <= "000000";
		when "000111000101010" => rgb <= "000000";
		when "000111000101110" => rgb <= "000000";
		when "000111000101111" => rgb <= "000000";
		when "000111000110000" => rgb <= "000000";
		when "000111000110001" => rgb <= "000000";
		when "000111000110010" => rgb <= "000000";
		when "000111000110011" => rgb <= "000000";
		when "000111000110111" => rgb <= "000000";
		when "000111000111000" => rgb <= "000000";
		when "000111000111001" => rgb <= "000000";
		when "000111000111010" => rgb <= "000000";
		when "000111000111011" => rgb <= "000000";
		when "000111000111100" => rgb <= "000000";
		when "000111000111101" => rgb <= "000000";
		when "000111000111110" => rgb <= "000000";
		when "000111000111111" => rgb <= "000000";
		when "000111001000000" => rgb <= "000000";
		when "000111001000001" => rgb <= "000000";
		when "000111001000010" => rgb <= "000000";
		when "000111001000011" => rgb <= "000000";
		when "000111001000100" => rgb <= "000000";
		when "000111001000101" => rgb <= "000000";
		when "000111001000110" => rgb <= "000000";
		when "000111001000111" => rgb <= "000000";
		when "000111001001000" => rgb <= "000000";
		when "000111001010110" => rgb <= "000000";
		when "000111001010111" => rgb <= "000000";
		when "000111001011000" => rgb <= "000000";
		when "000111001011001" => rgb <= "000000";
		when "000111001011010" => rgb <= "000000";
		when "000111001011011" => rgb <= "000000";
		when "000111001011100" => rgb <= "000000";
		when "000111001011101" => rgb <= "000000";
		when "000111001011110" => rgb <= "000000";
		when "000111001100010" => rgb <= "000000";
		when "000111001100011" => rgb <= "000000";
		when "000111001100100" => rgb <= "000000";
		when "000111001100101" => rgb <= "000000";
		when "000111001100110" => rgb <= "000000";
		when "000111001101011" => rgb <= "000000";
		when "000111001101100" => rgb <= "000000";
		when "000111001101101" => rgb <= "000000";
		when "000111001101110" => rgb <= "000000";
		when "000111001101111" => rgb <= "000000";
		when "000111001110001" => rgb <= "000000";
		when "000111001110010" => rgb <= "000000";
		when "000111001110011" => rgb <= "000000";
		when "000111001110100" => rgb <= "000000";
		when "000111001110101" => rgb <= "000000";
		when "000111001110110" => rgb <= "000000";
		when "000111001110111" => rgb <= "000000";
		when "000111001111000" => rgb <= "000000";
		when "000111001111001" => rgb <= "000000";
		when "000111001111010" => rgb <= "000000";
		when "000111001111011" => rgb <= "000000";
		when "000111001111100" => rgb <= "000000";
		when "000111001111110" => rgb <= "000000";
		when "000111001111111" => rgb <= "000000";
		when "000111010000000" => rgb <= "000000";
		when "000111010000001" => rgb <= "000000";
		when "000111010000010" => rgb <= "000000";
		when "000111010000011" => rgb <= "000000";
		when "000111010000100" => rgb <= "000000";
		when "000111010000101" => rgb <= "000000";
		when "000111010000110" => rgb <= "000000";
		when "000111010000111" => rgb <= "000000";
		when "000111010001000" => rgb <= "000000";
		when "000111010001001" => rgb <= "000000";
		when "000111100010011" => rgb <= "000000";
		when "000111100010100" => rgb <= "000000";
		when "000111100010101" => rgb <= "000000";
		when "000111100010110" => rgb <= "100110";
		when "000111100010111" => rgb <= "100110";
		when "000111100011000" => rgb <= "100110";
		when "000111100011001" => rgb <= "100110";
		when "000111100011010" => rgb <= "100110";
		when "000111100011011" => rgb <= "100110";
		when "000111100011100" => rgb <= "100110";
		when "000111100011101" => rgb <= "100110";
		when "000111100011110" => rgb <= "000000";
		when "000111100011111" => rgb <= "000000";
		when "000111100100011" => rgb <= "000000";
		when "000111100100100" => rgb <= "100110";
		when "000111100100101" => rgb <= "100110";
		when "000111100100110" => rgb <= "100110";
		when "000111100100111" => rgb <= "100110";
		when "000111100101000" => rgb <= "100110";
		when "000111100101001" => rgb <= "100110";
		when "000111100101010" => rgb <= "000000";
		when "000111100101011" => rgb <= "000000";
		when "000111100101100" => rgb <= "000000";
		when "000111100101110" => rgb <= "000000";
		when "000111100101111" => rgb <= "100110";
		when "000111100110000" => rgb <= "100110";
		when "000111100110001" => rgb <= "100110";
		when "000111100110010" => rgb <= "100110";
		when "000111100110011" => rgb <= "000000";
		when "000111100110100" => rgb <= "000000";
		when "000111100110111" => rgb <= "000000";
		when "000111100111000" => rgb <= "100110";
		when "000111100111001" => rgb <= "100110";
		when "000111100111010" => rgb <= "100110";
		when "000111100111011" => rgb <= "100110";
		when "000111100111100" => rgb <= "000000";
		when "000111100111101" => rgb <= "000000";
		when "000111100111110" => rgb <= "100110";
		when "000111100111111" => rgb <= "100110";
		when "000111101000000" => rgb <= "100110";
		when "000111101000001" => rgb <= "100110";
		when "000111101000010" => rgb <= "100110";
		when "000111101000011" => rgb <= "100110";
		when "000111101000100" => rgb <= "100110";
		when "000111101000101" => rgb <= "100110";
		when "000111101000110" => rgb <= "100110";
		when "000111101000111" => rgb <= "100110";
		when "000111101001000" => rgb <= "000000";
		when "000111101001001" => rgb <= "000000";
		when "000111101001010" => rgb <= "000000";
		when "000111101010100" => rgb <= "000000";
		when "000111101010101" => rgb <= "000000";
		when "000111101010110" => rgb <= "000000";
		when "000111101010111" => rgb <= "100110";
		when "000111101011000" => rgb <= "100110";
		when "000111101011001" => rgb <= "100110";
		when "000111101011010" => rgb <= "100110";
		when "000111101011011" => rgb <= "100110";
		when "000111101011100" => rgb <= "100110";
		when "000111101011101" => rgb <= "000000";
		when "000111101011110" => rgb <= "000000";
		when "000111101011111" => rgb <= "000000";
		when "000111101100010" => rgb <= "000000";
		when "000111101100011" => rgb <= "100110";
		when "000111101100100" => rgb <= "100110";
		when "000111101100101" => rgb <= "100110";
		when "000111101100110" => rgb <= "000000";
		when "000111101100111" => rgb <= "000000";
		when "000111101101000" => rgb <= "000000";
		when "000111101101011" => rgb <= "000000";
		when "000111101101100" => rgb <= "100110";
		when "000111101101101" => rgb <= "100110";
		when "000111101101110" => rgb <= "100110";
		when "000111101101111" => rgb <= "000000";
		when "000111101110000" => rgb <= "000000";
		when "000111101110001" => rgb <= "000000";
		when "000111101110010" => rgb <= "100110";
		when "000111101110011" => rgb <= "100110";
		when "000111101110100" => rgb <= "100110";
		when "000111101110101" => rgb <= "100110";
		when "000111101110110" => rgb <= "100110";
		when "000111101110111" => rgb <= "100110";
		when "000111101111000" => rgb <= "100110";
		when "000111101111001" => rgb <= "100110";
		when "000111101111010" => rgb <= "100110";
		when "000111101111011" => rgb <= "100110";
		when "000111101111100" => rgb <= "000000";
		when "000111101111101" => rgb <= "000000";
		when "000111101111110" => rgb <= "000000";
		when "000111101111111" => rgb <= "100110";
		when "000111110000000" => rgb <= "100110";
		when "000111110000001" => rgb <= "100110";
		when "000111110000010" => rgb <= "100110";
		when "000111110000011" => rgb <= "100110";
		when "000111110000100" => rgb <= "100110";
		when "000111110000101" => rgb <= "100110";
		when "000111110000110" => rgb <= "100110";
		when "000111110000111" => rgb <= "100110";
		when "000111110001000" => rgb <= "000000";
		when "000111110001001" => rgb <= "000000";
		when "000111110001010" => rgb <= "000000";
		when "000111110001011" => rgb <= "000000";
		when "001000000010010" => rgb <= "000000";
		when "001000000010011" => rgb <= "000000";
		when "001000000010100" => rgb <= "100110";
		when "001000000010101" => rgb <= "100110";
		when "001000000010110" => rgb <= "100110";
		when "001000000010111" => rgb <= "100110";
		when "001000000011000" => rgb <= "100110";
		when "001000000011001" => rgb <= "100110";
		when "001000000011010" => rgb <= "100110";
		when "001000000011011" => rgb <= "100110";
		when "001000000011100" => rgb <= "100110";
		when "001000000011101" => rgb <= "100110";
		when "001000000011110" => rgb <= "100110";
		when "001000000011111" => rgb <= "000000";
		when "001000000100000" => rgb <= "000000";
		when "001000000100001" => rgb <= "000000";
		when "001000000100010" => rgb <= "000000";
		when "001000000100011" => rgb <= "000000";
		when "001000000100100" => rgb <= "100110";
		when "001000000100101" => rgb <= "100110";
		when "001000000100110" => rgb <= "100110";
		when "001000000100111" => rgb <= "100110";
		when "001000000101000" => rgb <= "100110";
		when "001000000101001" => rgb <= "100110";
		when "001000000101010" => rgb <= "000000";
		when "001000000101011" => rgb <= "000000";
		when "001000000101100" => rgb <= "000000";
		when "001000000101101" => rgb <= "000000";
		when "001000000101110" => rgb <= "000000";
		when "001000000101111" => rgb <= "100110";
		when "001000000110000" => rgb <= "100110";
		when "001000000110001" => rgb <= "100110";
		when "001000000110010" => rgb <= "100110";
		when "001000000110011" => rgb <= "000000";
		when "001000000110100" => rgb <= "000000";
		when "001000000110101" => rgb <= "000000";
		when "001000000110110" => rgb <= "000000";
		when "001000000110111" => rgb <= "000000";
		when "001000000111000" => rgb <= "100110";
		when "001000000111001" => rgb <= "100110";
		when "001000000111010" => rgb <= "100110";
		when "001000000111011" => rgb <= "100110";
		when "001000000111100" => rgb <= "000000";
		when "001000000111101" => rgb <= "000000";
		when "001000000111110" => rgb <= "100110";
		when "001000000111111" => rgb <= "100110";
		when "001000001000000" => rgb <= "100110";
		when "001000001000001" => rgb <= "100110";
		when "001000001000010" => rgb <= "100110";
		when "001000001000011" => rgb <= "100110";
		when "001000001000100" => rgb <= "100110";
		when "001000001000101" => rgb <= "100110";
		when "001000001000110" => rgb <= "100110";
		when "001000001000111" => rgb <= "100110";
		when "001000001001000" => rgb <= "000000";
		when "001000001001001" => rgb <= "000000";
		when "001000001001010" => rgb <= "000000";
		when "001000001010100" => rgb <= "000000";
		when "001000001010101" => rgb <= "100110";
		when "001000001010110" => rgb <= "100110";
		when "001000001010111" => rgb <= "100110";
		when "001000001011000" => rgb <= "100110";
		when "001000001011001" => rgb <= "100110";
		when "001000001011010" => rgb <= "100110";
		when "001000001011011" => rgb <= "100110";
		when "001000001011100" => rgb <= "100110";
		when "001000001011101" => rgb <= "100110";
		when "001000001011110" => rgb <= "100110";
		when "001000001011111" => rgb <= "000000";
		when "001000001100000" => rgb <= "000000";
		when "001000001100010" => rgb <= "000000";
		when "001000001100011" => rgb <= "100110";
		when "001000001100100" => rgb <= "100110";
		when "001000001100101" => rgb <= "100110";
		when "001000001100110" => rgb <= "000000";
		when "001000001100111" => rgb <= "000000";
		when "001000001101000" => rgb <= "000000";
		when "001000001101011" => rgb <= "000000";
		when "001000001101100" => rgb <= "100110";
		when "001000001101101" => rgb <= "100110";
		when "001000001101110" => rgb <= "100110";
		when "001000001101111" => rgb <= "000000";
		when "001000001110000" => rgb <= "000000";
		when "001000001110001" => rgb <= "000000";
		when "001000001110010" => rgb <= "100110";
		when "001000001110011" => rgb <= "100110";
		when "001000001110100" => rgb <= "100110";
		when "001000001110101" => rgb <= "100110";
		when "001000001110110" => rgb <= "100110";
		when "001000001110111" => rgb <= "100110";
		when "001000001111000" => rgb <= "100110";
		when "001000001111001" => rgb <= "100110";
		when "001000001111010" => rgb <= "100110";
		when "001000001111011" => rgb <= "100110";
		when "001000001111100" => rgb <= "000000";
		when "001000001111101" => rgb <= "000000";
		when "001000001111110" => rgb <= "000000";
		when "001000001111111" => rgb <= "100110";
		when "001000010000000" => rgb <= "100110";
		when "001000010000001" => rgb <= "100110";
		when "001000010000010" => rgb <= "100110";
		when "001000010000011" => rgb <= "100110";
		when "001000010000100" => rgb <= "100110";
		when "001000010000101" => rgb <= "100110";
		when "001000010000110" => rgb <= "100110";
		when "001000010000111" => rgb <= "100110";
		when "001000010001000" => rgb <= "100110";
		when "001000010001001" => rgb <= "100110";
		when "001000010001010" => rgb <= "000000";
		when "001000010001011" => rgb <= "000000";
		when "001000010001100" => rgb <= "000000";
		when "001000100010010" => rgb <= "000000";
		when "001000100010011" => rgb <= "100110";
		when "001000100010100" => rgb <= "100110";
		when "001000100010101" => rgb <= "100110";
		when "001000100010110" => rgb <= "100110";
		when "001000100010111" => rgb <= "100110";
		when "001000100011000" => rgb <= "100110";
		when "001000100011001" => rgb <= "100110";
		when "001000100011010" => rgb <= "100110";
		when "001000100011011" => rgb <= "100110";
		when "001000100011100" => rgb <= "100110";
		when "001000100011101" => rgb <= "100110";
		when "001000100011110" => rgb <= "100110";
		when "001000100011111" => rgb <= "000000";
		when "001000100100000" => rgb <= "000000";
		when "001000100100001" => rgb <= "000000";
		when "001000100100010" => rgb <= "100110";
		when "001000100100011" => rgb <= "100110";
		when "001000100100100" => rgb <= "100110";
		when "001000100100101" => rgb <= "100110";
		when "001000100100110" => rgb <= "100110";
		when "001000100100111" => rgb <= "100110";
		when "001000100101000" => rgb <= "100110";
		when "001000100101001" => rgb <= "100110";
		when "001000100101010" => rgb <= "100110";
		when "001000100101011" => rgb <= "100110";
		when "001000100101100" => rgb <= "000000";
		when "001000100101101" => rgb <= "000000";
		when "001000100101110" => rgb <= "000000";
		when "001000100101111" => rgb <= "100110";
		when "001000100110000" => rgb <= "100110";
		when "001000100110001" => rgb <= "100110";
		when "001000100110010" => rgb <= "100110";
		when "001000100110011" => rgb <= "100110";
		when "001000100110100" => rgb <= "000000";
		when "001000100110101" => rgb <= "000000";
		when "001000100110110" => rgb <= "000000";
		when "001000100110111" => rgb <= "100110";
		when "001000100111000" => rgb <= "100110";
		when "001000100111001" => rgb <= "100110";
		when "001000100111010" => rgb <= "100110";
		when "001000100111011" => rgb <= "100110";
		when "001000100111100" => rgb <= "000000";
		when "001000100111101" => rgb <= "000000";
		when "001000100111110" => rgb <= "100110";
		when "001000100111111" => rgb <= "100110";
		when "001000101000000" => rgb <= "100110";
		when "001000101000001" => rgb <= "100110";
		when "001000101000010" => rgb <= "100110";
		when "001000101000011" => rgb <= "100110";
		when "001000101000100" => rgb <= "100110";
		when "001000101000101" => rgb <= "100110";
		when "001000101000110" => rgb <= "100110";
		when "001000101000111" => rgb <= "100110";
		when "001000101001000" => rgb <= "000000";
		when "001000101001001" => rgb <= "000000";
		when "001000101001010" => rgb <= "000000";
		when "001000101010011" => rgb <= "000000";
		when "001000101010100" => rgb <= "000000";
		when "001000101010101" => rgb <= "100110";
		when "001000101010110" => rgb <= "100110";
		when "001000101010111" => rgb <= "100110";
		when "001000101011000" => rgb <= "100110";
		when "001000101011001" => rgb <= "100110";
		when "001000101011010" => rgb <= "100110";
		when "001000101011011" => rgb <= "100110";
		when "001000101011100" => rgb <= "100110";
		when "001000101011101" => rgb <= "100110";
		when "001000101011110" => rgb <= "100110";
		when "001000101011111" => rgb <= "000000";
		when "001000101100000" => rgb <= "000000";
		when "001000101100001" => rgb <= "000000";
		when "001000101100010" => rgb <= "000000";
		when "001000101100011" => rgb <= "100110";
		when "001000101100100" => rgb <= "100110";
		when "001000101100101" => rgb <= "100110";
		when "001000101100110" => rgb <= "000000";
		when "001000101100111" => rgb <= "000000";
		when "001000101101000" => rgb <= "000000";
		when "001000101101011" => rgb <= "000000";
		when "001000101101100" => rgb <= "100110";
		when "001000101101101" => rgb <= "100110";
		when "001000101101110" => rgb <= "100110";
		when "001000101101111" => rgb <= "000000";
		when "001000101110000" => rgb <= "000000";
		when "001000101110001" => rgb <= "000000";
		when "001000101110010" => rgb <= "100110";
		when "001000101110011" => rgb <= "100110";
		when "001000101110100" => rgb <= "100110";
		when "001000101110101" => rgb <= "100110";
		when "001000101110110" => rgb <= "100110";
		when "001000101110111" => rgb <= "100110";
		when "001000101111000" => rgb <= "100110";
		when "001000101111001" => rgb <= "100110";
		when "001000101111010" => rgb <= "100110";
		when "001000101111011" => rgb <= "100110";
		when "001000101111100" => rgb <= "000000";
		when "001000101111101" => rgb <= "000000";
		when "001000101111110" => rgb <= "000000";
		when "001000101111111" => rgb <= "100110";
		when "001000110000000" => rgb <= "100110";
		when "001000110000001" => rgb <= "100110";
		when "001000110000010" => rgb <= "000000";
		when "001000110000011" => rgb <= "000000";
		when "001000110000100" => rgb <= "000000";
		when "001000110000101" => rgb <= "000000";
		when "001000110000110" => rgb <= "000000";
		when "001000110000111" => rgb <= "100110";
		when "001000110001000" => rgb <= "100110";
		when "001000110001001" => rgb <= "100110";
		when "001000110001010" => rgb <= "000000";
		when "001000110001011" => rgb <= "000000";
		when "001000110001100" => rgb <= "000000";
		when "001001000010010" => rgb <= "000000";
		when "001001000010011" => rgb <= "100110";
		when "001001000010100" => rgb <= "100110";
		when "001001000010101" => rgb <= "100110";
		when "001001000010110" => rgb <= "100110";
		when "001001000010111" => rgb <= "000000";
		when "001001000011000" => rgb <= "000000";
		when "001001000011001" => rgb <= "000000";
		when "001001000011010" => rgb <= "000000";
		when "001001000011011" => rgb <= "000000";
		when "001001000011100" => rgb <= "100110";
		when "001001000011101" => rgb <= "100110";
		when "001001000011110" => rgb <= "100110";
		when "001001000011111" => rgb <= "000000";
		when "001001000100000" => rgb <= "000000";
		when "001001000100001" => rgb <= "000000";
		when "001001000100010" => rgb <= "100110";
		when "001001000100011" => rgb <= "100110";
		when "001001000100100" => rgb <= "100110";
		when "001001000100101" => rgb <= "000000";
		when "001001000100110" => rgb <= "000000";
		when "001001000100111" => rgb <= "000000";
		when "001001000101000" => rgb <= "000000";
		when "001001000101001" => rgb <= "100110";
		when "001001000101010" => rgb <= "100110";
		when "001001000101011" => rgb <= "100110";
		when "001001000101100" => rgb <= "000000";
		when "001001000101101" => rgb <= "000000";
		when "001001000101110" => rgb <= "000000";
		when "001001000101111" => rgb <= "100110";
		when "001001000110000" => rgb <= "100110";
		when "001001000110001" => rgb <= "100110";
		when "001001000110010" => rgb <= "100110";
		when "001001000110011" => rgb <= "100110";
		when "001001000110100" => rgb <= "000000";
		when "001001000110101" => rgb <= "000000";
		when "001001000110110" => rgb <= "000000";
		when "001001000110111" => rgb <= "100110";
		when "001001000111000" => rgb <= "100110";
		when "001001000111001" => rgb <= "100110";
		when "001001000111010" => rgb <= "100110";
		when "001001000111011" => rgb <= "100110";
		when "001001000111100" => rgb <= "000000";
		when "001001000111101" => rgb <= "000000";
		when "001001000111110" => rgb <= "100110";
		when "001001000111111" => rgb <= "100110";
		when "001001001000000" => rgb <= "100110";
		when "001001001000001" => rgb <= "000000";
		when "001001001000010" => rgb <= "000000";
		when "001001001000011" => rgb <= "000000";
		when "001001001000100" => rgb <= "000000";
		when "001001001000101" => rgb <= "000000";
		when "001001001000110" => rgb <= "000000";
		when "001001001000111" => rgb <= "000000";
		when "001001001001000" => rgb <= "000000";
		when "001001001001001" => rgb <= "000000";
		when "001001001001010" => rgb <= "000000";
		when "001001001010011" => rgb <= "000000";
		when "001001001010100" => rgb <= "100110";
		when "001001001010101" => rgb <= "100110";
		when "001001001010110" => rgb <= "100110";
		when "001001001010111" => rgb <= "100110";
		when "001001001011000" => rgb <= "000000";
		when "001001001011001" => rgb <= "000000";
		when "001001001011010" => rgb <= "000000";
		when "001001001011011" => rgb <= "000000";
		when "001001001011100" => rgb <= "100110";
		when "001001001011101" => rgb <= "100110";
		when "001001001011110" => rgb <= "100110";
		when "001001001011111" => rgb <= "100110";
		when "001001001100000" => rgb <= "000000";
		when "001001001100001" => rgb <= "000000";
		when "001001001100010" => rgb <= "000000";
		when "001001001100011" => rgb <= "100110";
		when "001001001100100" => rgb <= "100110";
		when "001001001100101" => rgb <= "100110";
		when "001001001100110" => rgb <= "000000";
		when "001001001100111" => rgb <= "000000";
		when "001001001101000" => rgb <= "000000";
		when "001001001101011" => rgb <= "000000";
		when "001001001101100" => rgb <= "100110";
		when "001001001101101" => rgb <= "100110";
		when "001001001101110" => rgb <= "100110";
		when "001001001101111" => rgb <= "000000";
		when "001001001110000" => rgb <= "000000";
		when "001001001110001" => rgb <= "000000";
		when "001001001110010" => rgb <= "100110";
		when "001001001110011" => rgb <= "100110";
		when "001001001110100" => rgb <= "100110";
		when "001001001110101" => rgb <= "000000";
		when "001001001110110" => rgb <= "000000";
		when "001001001110111" => rgb <= "000000";
		when "001001001111000" => rgb <= "000000";
		when "001001001111001" => rgb <= "000000";
		when "001001001111010" => rgb <= "000000";
		when "001001001111011" => rgb <= "000000";
		when "001001001111100" => rgb <= "000000";
		when "001001001111101" => rgb <= "000000";
		when "001001001111110" => rgb <= "000000";
		when "001001001111111" => rgb <= "100110";
		when "001001010000000" => rgb <= "100110";
		when "001001010000001" => rgb <= "100110";
		when "001001010000010" => rgb <= "000000";
		when "001001010000011" => rgb <= "000000";
		when "001001010000100" => rgb <= "000000";
		when "001001010000101" => rgb <= "000000";
		when "001001010000110" => rgb <= "000000";
		when "001001010000111" => rgb <= "100110";
		when "001001010001000" => rgb <= "100110";
		when "001001010001001" => rgb <= "100110";
		when "001001010001010" => rgb <= "000000";
		when "001001010001011" => rgb <= "000000";
		when "001001010001100" => rgb <= "000000";
		when "001001100010010" => rgb <= "000000";
		when "001001100010011" => rgb <= "100110";
		when "001001100010100" => rgb <= "100110";
		when "001001100010101" => rgb <= "100110";
		when "001001100010110" => rgb <= "000000";
		when "001001100010111" => rgb <= "000000";
		when "001001100011000" => rgb <= "000000";
		when "001001100011001" => rgb <= "000000";
		when "001001100011010" => rgb <= "000000";
		when "001001100011011" => rgb <= "000000";
		when "001001100011100" => rgb <= "000000";
		when "001001100011101" => rgb <= "000000";
		when "001001100011110" => rgb <= "000000";
		when "001001100011111" => rgb <= "000000";
		when "001001100100000" => rgb <= "000000";
		when "001001100100001" => rgb <= "000000";
		when "001001100100010" => rgb <= "100110";
		when "001001100100011" => rgb <= "100110";
		when "001001100100100" => rgb <= "100110";
		when "001001100100101" => rgb <= "000000";
		when "001001100100110" => rgb <= "000000";
		when "001001100100111" => rgb <= "000000";
		when "001001100101000" => rgb <= "000000";
		when "001001100101001" => rgb <= "100110";
		when "001001100101010" => rgb <= "100110";
		when "001001100101011" => rgb <= "100110";
		when "001001100101100" => rgb <= "000000";
		when "001001100101101" => rgb <= "000000";
		when "001001100101110" => rgb <= "000000";
		when "001001100101111" => rgb <= "100110";
		when "001001100110000" => rgb <= "100110";
		when "001001100110001" => rgb <= "100110";
		when "001001100110010" => rgb <= "100110";
		when "001001100110011" => rgb <= "100110";
		when "001001100110100" => rgb <= "100110";
		when "001001100110101" => rgb <= "000000";
		when "001001100110110" => rgb <= "100110";
		when "001001100110111" => rgb <= "100110";
		when "001001100111000" => rgb <= "100110";
		when "001001100111001" => rgb <= "100110";
		when "001001100111010" => rgb <= "100110";
		when "001001100111011" => rgb <= "100110";
		when "001001100111100" => rgb <= "000000";
		when "001001100111101" => rgb <= "000000";
		when "001001100111110" => rgb <= "100110";
		when "001001100111111" => rgb <= "100110";
		when "001001101000000" => rgb <= "100110";
		when "001001101000001" => rgb <= "000000";
		when "001001101000010" => rgb <= "000000";
		when "001001101000011" => rgb <= "000000";
		when "001001101000100" => rgb <= "000000";
		when "001001101000101" => rgb <= "000000";
		when "001001101000110" => rgb <= "000000";
		when "001001101000111" => rgb <= "000000";
		when "001001101001000" => rgb <= "000000";
		when "001001101001001" => rgb <= "000000";
		when "001001101001010" => rgb <= "000000";
		when "001001101010011" => rgb <= "000000";
		when "001001101010100" => rgb <= "100110";
		when "001001101010101" => rgb <= "100110";
		when "001001101010110" => rgb <= "100110";
		when "001001101010111" => rgb <= "000000";
		when "001001101011000" => rgb <= "000000";
		when "001001101011001" => rgb <= "000000";
		when "001001101011010" => rgb <= "000000";
		when "001001101011011" => rgb <= "000000";
		when "001001101011100" => rgb <= "000000";
		when "001001101011101" => rgb <= "100110";
		when "001001101011110" => rgb <= "100110";
		when "001001101011111" => rgb <= "100110";
		when "001001101100000" => rgb <= "000000";
		when "001001101100001" => rgb <= "000000";
		when "001001101100010" => rgb <= "000000";
		when "001001101100011" => rgb <= "100110";
		when "001001101100100" => rgb <= "100110";
		when "001001101100101" => rgb <= "100110";
		when "001001101100110" => rgb <= "000000";
		when "001001101100111" => rgb <= "000000";
		when "001001101101000" => rgb <= "000000";
		when "001001101101011" => rgb <= "000000";
		when "001001101101100" => rgb <= "100110";
		when "001001101101101" => rgb <= "100110";
		when "001001101101110" => rgb <= "100110";
		when "001001101101111" => rgb <= "000000";
		when "001001101110000" => rgb <= "000000";
		when "001001101110001" => rgb <= "000000";
		when "001001101110010" => rgb <= "100110";
		when "001001101110011" => rgb <= "100110";
		when "001001101110100" => rgb <= "100110";
		when "001001101110101" => rgb <= "000000";
		when "001001101110110" => rgb <= "000000";
		when "001001101110111" => rgb <= "000000";
		when "001001101111000" => rgb <= "000000";
		when "001001101111001" => rgb <= "000000";
		when "001001101111010" => rgb <= "000000";
		when "001001101111011" => rgb <= "000000";
		when "001001101111100" => rgb <= "000000";
		when "001001101111101" => rgb <= "000000";
		when "001001101111110" => rgb <= "000000";
		when "001001101111111" => rgb <= "100110";
		when "001001110000000" => rgb <= "100110";
		when "001001110000001" => rgb <= "100110";
		when "001001110000010" => rgb <= "000000";
		when "001001110000011" => rgb <= "000000";
		when "001001110000100" => rgb <= "000000";
		when "001001110000101" => rgb <= "000000";
		when "001001110000110" => rgb <= "000000";
		when "001001110000111" => rgb <= "100110";
		when "001001110001000" => rgb <= "100110";
		when "001001110001001" => rgb <= "100110";
		when "001001110001010" => rgb <= "000000";
		when "001001110001011" => rgb <= "000000";
		when "001001110001100" => rgb <= "000000";
		when "001010000010010" => rgb <= "000000";
		when "001010000010011" => rgb <= "100110";
		when "001010000010100" => rgb <= "100110";
		when "001010000010101" => rgb <= "100110";
		when "001010000010110" => rgb <= "000000";
		when "001010000010111" => rgb <= "000000";
		when "001010000011000" => rgb <= "000000";
		when "001010000011001" => rgb <= "000000";
		when "001010000011010" => rgb <= "000000";
		when "001010000011011" => rgb <= "000000";
		when "001010000011100" => rgb <= "000000";
		when "001010000011101" => rgb <= "000000";
		when "001010000011110" => rgb <= "000000";
		when "001010000011111" => rgb <= "000000";
		when "001010000100000" => rgb <= "000000";
		when "001010000100001" => rgb <= "100110";
		when "001010000100010" => rgb <= "100110";
		when "001010000100011" => rgb <= "100110";
		when "001010000100100" => rgb <= "000000";
		when "001010000100101" => rgb <= "000000";
		when "001010000100110" => rgb <= "000000";
		when "001010000100111" => rgb <= "000000";
		when "001010000101000" => rgb <= "000000";
		when "001010000101001" => rgb <= "000000";
		when "001010000101010" => rgb <= "100110";
		when "001010000101011" => rgb <= "100110";
		when "001010000101100" => rgb <= "100110";
		when "001010000101101" => rgb <= "000000";
		when "001010000101110" => rgb <= "000000";
		when "001010000101111" => rgb <= "100110";
		when "001010000110000" => rgb <= "100110";
		when "001010000110001" => rgb <= "100110";
		when "001010000110010" => rgb <= "100110";
		when "001010000110011" => rgb <= "100110";
		when "001010000110100" => rgb <= "100110";
		when "001010000110101" => rgb <= "100110";
		when "001010000110110" => rgb <= "100110";
		when "001010000110111" => rgb <= "100110";
		when "001010000111000" => rgb <= "100110";
		when "001010000111001" => rgb <= "100110";
		when "001010000111010" => rgb <= "100110";
		when "001010000111011" => rgb <= "100110";
		when "001010000111100" => rgb <= "000000";
		when "001010000111101" => rgb <= "000000";
		when "001010000111110" => rgb <= "100110";
		when "001010000111111" => rgb <= "100110";
		when "001010001000000" => rgb <= "100110";
		when "001010001000001" => rgb <= "000000";
		when "001010001000010" => rgb <= "000000";
		when "001010001000011" => rgb <= "000000";
		when "001010001000100" => rgb <= "000000";
		when "001010001000101" => rgb <= "000000";
		when "001010001000110" => rgb <= "000000";
		when "001010001000111" => rgb <= "000000";
		when "001010001001000" => rgb <= "000000";
		when "001010001010011" => rgb <= "000000";
		when "001010001010100" => rgb <= "100110";
		when "001010001010101" => rgb <= "100110";
		when "001010001010110" => rgb <= "100110";
		when "001010001010111" => rgb <= "000000";
		when "001010001011000" => rgb <= "000000";
		when "001010001011001" => rgb <= "000000";
		when "001010001011010" => rgb <= "000000";
		when "001010001011011" => rgb <= "000000";
		when "001010001011100" => rgb <= "000000";
		when "001010001011101" => rgb <= "100110";
		when "001010001011110" => rgb <= "100110";
		when "001010001011111" => rgb <= "100110";
		when "001010001100000" => rgb <= "000000";
		when "001010001100001" => rgb <= "000000";
		when "001010001100010" => rgb <= "000000";
		when "001010001100011" => rgb <= "100110";
		when "001010001100100" => rgb <= "100110";
		when "001010001100101" => rgb <= "100110";
		when "001010001100110" => rgb <= "000000";
		when "001010001100111" => rgb <= "000000";
		when "001010001101000" => rgb <= "000000";
		when "001010001101011" => rgb <= "000000";
		when "001010001101100" => rgb <= "100110";
		when "001010001101101" => rgb <= "100110";
		when "001010001101110" => rgb <= "100110";
		when "001010001101111" => rgb <= "000000";
		when "001010001110000" => rgb <= "000000";
		when "001010001110001" => rgb <= "000000";
		when "001010001110010" => rgb <= "100110";
		when "001010001110011" => rgb <= "100110";
		when "001010001110100" => rgb <= "100110";
		when "001010001110101" => rgb <= "000000";
		when "001010001110110" => rgb <= "000000";
		when "001010001110111" => rgb <= "000000";
		when "001010001111000" => rgb <= "000000";
		when "001010001111001" => rgb <= "000000";
		when "001010001111010" => rgb <= "000000";
		when "001010001111011" => rgb <= "000000";
		when "001010001111100" => rgb <= "000000";
		when "001010001111110" => rgb <= "000000";
		when "001010001111111" => rgb <= "100110";
		when "001010010000000" => rgb <= "100110";
		when "001010010000001" => rgb <= "100110";
		when "001010010000010" => rgb <= "000000";
		when "001010010000011" => rgb <= "000000";
		when "001010010000100" => rgb <= "000000";
		when "001010010000101" => rgb <= "000000";
		when "001010010000110" => rgb <= "000000";
		when "001010010000111" => rgb <= "100110";
		when "001010010001000" => rgb <= "100110";
		when "001010010001001" => rgb <= "100110";
		when "001010010001010" => rgb <= "000000";
		when "001010010001011" => rgb <= "000000";
		when "001010010001100" => rgb <= "000000";
		when "001010100010010" => rgb <= "000000";
		when "001010100010011" => rgb <= "100110";
		when "001010100010100" => rgb <= "100110";
		when "001010100010101" => rgb <= "100110";
		when "001010100010110" => rgb <= "000000";
		when "001010100010111" => rgb <= "000000";
		when "001010100011000" => rgb <= "000000";
		when "001010100011001" => rgb <= "100110";
		when "001010100011010" => rgb <= "100110";
		when "001010100011011" => rgb <= "100110";
		when "001010100011100" => rgb <= "100110";
		when "001010100011101" => rgb <= "100110";
		when "001010100011110" => rgb <= "100110";
		when "001010100011111" => rgb <= "000000";
		when "001010100100000" => rgb <= "000000";
		when "001010100100001" => rgb <= "100110";
		when "001010100100010" => rgb <= "100110";
		when "001010100100011" => rgb <= "100110";
		when "001010100100100" => rgb <= "000000";
		when "001010100100101" => rgb <= "000000";
		when "001010100100110" => rgb <= "000000";
		when "001010100100111" => rgb <= "000000";
		when "001010100101000" => rgb <= "000000";
		when "001010100101001" => rgb <= "000000";
		when "001010100101010" => rgb <= "100110";
		when "001010100101011" => rgb <= "100110";
		when "001010100101100" => rgb <= "100110";
		when "001010100101101" => rgb <= "000000";
		when "001010100101110" => rgb <= "000000";
		when "001010100101111" => rgb <= "100110";
		when "001010100110000" => rgb <= "100110";
		when "001010100110001" => rgb <= "100110";
		when "001010100110010" => rgb <= "000000";
		when "001010100110011" => rgb <= "100110";
		when "001010100110100" => rgb <= "100110";
		when "001010100110101" => rgb <= "100110";
		when "001010100110110" => rgb <= "100110";
		when "001010100110111" => rgb <= "100110";
		when "001010100111000" => rgb <= "000000";
		when "001010100111001" => rgb <= "100110";
		when "001010100111010" => rgb <= "100110";
		when "001010100111011" => rgb <= "100110";
		when "001010100111100" => rgb <= "000000";
		when "001010100111101" => rgb <= "000000";
		when "001010100111110" => rgb <= "100110";
		when "001010100111111" => rgb <= "100110";
		when "001010101000000" => rgb <= "100110";
		when "001010101000001" => rgb <= "100110";
		when "001010101000010" => rgb <= "100110";
		when "001010101000011" => rgb <= "100110";
		when "001010101000100" => rgb <= "100110";
		when "001010101000101" => rgb <= "100110";
		when "001010101000110" => rgb <= "100110";
		when "001010101000111" => rgb <= "000000";
		when "001010101001000" => rgb <= "000000";
		when "001010101010011" => rgb <= "000000";
		when "001010101010100" => rgb <= "100110";
		when "001010101010101" => rgb <= "100110";
		when "001010101010110" => rgb <= "100110";
		when "001010101010111" => rgb <= "000000";
		when "001010101011000" => rgb <= "000000";
		when "001010101011001" => rgb <= "000000";
		when "001010101011010" => rgb <= "000000";
		when "001010101011011" => rgb <= "000000";
		when "001010101011100" => rgb <= "000000";
		when "001010101011101" => rgb <= "100110";
		when "001010101011110" => rgb <= "100110";
		when "001010101011111" => rgb <= "100110";
		when "001010101100000" => rgb <= "000000";
		when "001010101100001" => rgb <= "000000";
		when "001010101100010" => rgb <= "000000";
		when "001010101100011" => rgb <= "100110";
		when "001010101100100" => rgb <= "100110";
		when "001010101100101" => rgb <= "100110";
		when "001010101100110" => rgb <= "000000";
		when "001010101100111" => rgb <= "000000";
		when "001010101101000" => rgb <= "000000";
		when "001010101101001" => rgb <= "000000";
		when "001010101101011" => rgb <= "000000";
		when "001010101101100" => rgb <= "100110";
		when "001010101101101" => rgb <= "100110";
		when "001010101101110" => rgb <= "100110";
		when "001010101101111" => rgb <= "000000";
		when "001010101110000" => rgb <= "000000";
		when "001010101110001" => rgb <= "000000";
		when "001010101110010" => rgb <= "100110";
		when "001010101110011" => rgb <= "100110";
		when "001010101110100" => rgb <= "100110";
		when "001010101110101" => rgb <= "100110";
		when "001010101110110" => rgb <= "100110";
		when "001010101110111" => rgb <= "100110";
		when "001010101111000" => rgb <= "100110";
		when "001010101111001" => rgb <= "100110";
		when "001010101111010" => rgb <= "100110";
		when "001010101111011" => rgb <= "000000";
		when "001010101111100" => rgb <= "000000";
		when "001010101111110" => rgb <= "000000";
		when "001010101111111" => rgb <= "100110";
		when "001010110000000" => rgb <= "100110";
		when "001010110000001" => rgb <= "100110";
		when "001010110000010" => rgb <= "000000";
		when "001010110000011" => rgb <= "000000";
		when "001010110000100" => rgb <= "000000";
		when "001010110000101" => rgb <= "000000";
		when "001010110000110" => rgb <= "100110";
		when "001010110000111" => rgb <= "100110";
		when "001010110001000" => rgb <= "100110";
		when "001010110001001" => rgb <= "100110";
		when "001010110001010" => rgb <= "000000";
		when "001010110001011" => rgb <= "000000";
		when "001010110001100" => rgb <= "000000";
		when "001011000010010" => rgb <= "000000";
		when "001011000010011" => rgb <= "100110";
		when "001011000010100" => rgb <= "100110";
		when "001011000010101" => rgb <= "100110";
		when "001011000010110" => rgb <= "000000";
		when "001011000010111" => rgb <= "000000";
		when "001011000011000" => rgb <= "000000";
		when "001011000011001" => rgb <= "100110";
		when "001011000011010" => rgb <= "100110";
		when "001011000011011" => rgb <= "100110";
		when "001011000011100" => rgb <= "100110";
		when "001011000011101" => rgb <= "100110";
		when "001011000011110" => rgb <= "100110";
		when "001011000011111" => rgb <= "000000";
		when "001011000100000" => rgb <= "000000";
		when "001011000100001" => rgb <= "100110";
		when "001011000100010" => rgb <= "100110";
		when "001011000100011" => rgb <= "100110";
		when "001011000100100" => rgb <= "100110";
		when "001011000100101" => rgb <= "100110";
		when "001011000100110" => rgb <= "100110";
		when "001011000100111" => rgb <= "100110";
		when "001011000101000" => rgb <= "100110";
		when "001011000101001" => rgb <= "100110";
		when "001011000101010" => rgb <= "100110";
		when "001011000101011" => rgb <= "100110";
		when "001011000101100" => rgb <= "100110";
		when "001011000101101" => rgb <= "000000";
		when "001011000101110" => rgb <= "000000";
		when "001011000101111" => rgb <= "100110";
		when "001011000110000" => rgb <= "100110";
		when "001011000110001" => rgb <= "100110";
		when "001011000110010" => rgb <= "000000";
		when "001011000110011" => rgb <= "100110";
		when "001011000110100" => rgb <= "100110";
		when "001011000110101" => rgb <= "100110";
		when "001011000110110" => rgb <= "100110";
		when "001011000110111" => rgb <= "100110";
		when "001011000111000" => rgb <= "000000";
		when "001011000111001" => rgb <= "100110";
		when "001011000111010" => rgb <= "100110";
		when "001011000111011" => rgb <= "100110";
		when "001011000111100" => rgb <= "000000";
		when "001011000111101" => rgb <= "000000";
		when "001011000111110" => rgb <= "100110";
		when "001011000111111" => rgb <= "100110";
		when "001011001000000" => rgb <= "100110";
		when "001011001000001" => rgb <= "100110";
		when "001011001000010" => rgb <= "100110";
		when "001011001000011" => rgb <= "100110";
		when "001011001000100" => rgb <= "100110";
		when "001011001000101" => rgb <= "100110";
		when "001011001000110" => rgb <= "100110";
		when "001011001000111" => rgb <= "000000";
		when "001011001001000" => rgb <= "000000";
		when "001011001010011" => rgb <= "000000";
		when "001011001010100" => rgb <= "100110";
		when "001011001010101" => rgb <= "100110";
		when "001011001010110" => rgb <= "100110";
		when "001011001010111" => rgb <= "000000";
		when "001011001011000" => rgb <= "000000";
		when "001011001011001" => rgb <= "000000";
		when "001011001011010" => rgb <= "000000";
		when "001011001011011" => rgb <= "000000";
		when "001011001011100" => rgb <= "000000";
		when "001011001011101" => rgb <= "100110";
		when "001011001011110" => rgb <= "100110";
		when "001011001011111" => rgb <= "100110";
		when "001011001100000" => rgb <= "000000";
		when "001011001100001" => rgb <= "000000";
		when "001011001100010" => rgb <= "000000";
		when "001011001100011" => rgb <= "000000";
		when "001011001100100" => rgb <= "100110";
		when "001011001100101" => rgb <= "100110";
		when "001011001100110" => rgb <= "000000";
		when "001011001100111" => rgb <= "000000";
		when "001011001101000" => rgb <= "000000";
		when "001011001101001" => rgb <= "000000";
		when "001011001101010" => rgb <= "000000";
		when "001011001101011" => rgb <= "000000";
		when "001011001101100" => rgb <= "100110";
		when "001011001101101" => rgb <= "100110";
		when "001011001101110" => rgb <= "000000";
		when "001011001101111" => rgb <= "000000";
		when "001011001110000" => rgb <= "000000";
		when "001011001110001" => rgb <= "000000";
		when "001011001110010" => rgb <= "100110";
		when "001011001110011" => rgb <= "100110";
		when "001011001110100" => rgb <= "100110";
		when "001011001110101" => rgb <= "100110";
		when "001011001110110" => rgb <= "100110";
		when "001011001110111" => rgb <= "100110";
		when "001011001111000" => rgb <= "100110";
		when "001011001111001" => rgb <= "100110";
		when "001011001111010" => rgb <= "100110";
		when "001011001111011" => rgb <= "000000";
		when "001011001111100" => rgb <= "000000";
		when "001011001111110" => rgb <= "000000";
		when "001011001111111" => rgb <= "100110";
		when "001011010000000" => rgb <= "100110";
		when "001011010000001" => rgb <= "100110";
		when "001011010000010" => rgb <= "100110";
		when "001011010000011" => rgb <= "100110";
		when "001011010000100" => rgb <= "100110";
		when "001011010000101" => rgb <= "100110";
		when "001011010000110" => rgb <= "100110";
		when "001011010000111" => rgb <= "100110";
		when "001011010001000" => rgb <= "000000";
		when "001011010001001" => rgb <= "000000";
		when "001011010001010" => rgb <= "000000";
		when "001011010001011" => rgb <= "000000";
		when "001011100010010" => rgb <= "000000";
		when "001011100010011" => rgb <= "100110";
		when "001011100010100" => rgb <= "100110";
		when "001011100010101" => rgb <= "100110";
		when "001011100010110" => rgb <= "000000";
		when "001011100010111" => rgb <= "000000";
		when "001011100011000" => rgb <= "000000";
		when "001011100011001" => rgb <= "000000";
		when "001011100011010" => rgb <= "000000";
		when "001011100011011" => rgb <= "000000";
		when "001011100011100" => rgb <= "100110";
		when "001011100011101" => rgb <= "100110";
		when "001011100011110" => rgb <= "100110";
		when "001011100011111" => rgb <= "000000";
		when "001011100100000" => rgb <= "000000";
		when "001011100100001" => rgb <= "100110";
		when "001011100100010" => rgb <= "100110";
		when "001011100100011" => rgb <= "100110";
		when "001011100100100" => rgb <= "100110";
		when "001011100100101" => rgb <= "100110";
		when "001011100100110" => rgb <= "100110";
		when "001011100100111" => rgb <= "100110";
		when "001011100101000" => rgb <= "100110";
		when "001011100101001" => rgb <= "100110";
		when "001011100101010" => rgb <= "100110";
		when "001011100101011" => rgb <= "100110";
		when "001011100101100" => rgb <= "100110";
		when "001011100101101" => rgb <= "000000";
		when "001011100101110" => rgb <= "000000";
		when "001011100101111" => rgb <= "100110";
		when "001011100110000" => rgb <= "100110";
		when "001011100110001" => rgb <= "100110";
		when "001011100110010" => rgb <= "000000";
		when "001011100110011" => rgb <= "000000";
		when "001011100110100" => rgb <= "100110";
		when "001011100110101" => rgb <= "100110";
		when "001011100110110" => rgb <= "100110";
		when "001011100110111" => rgb <= "000000";
		when "001011100111000" => rgb <= "000000";
		when "001011100111001" => rgb <= "100110";
		when "001011100111010" => rgb <= "100110";
		when "001011100111011" => rgb <= "100110";
		when "001011100111100" => rgb <= "000000";
		when "001011100111101" => rgb <= "000000";
		when "001011100111110" => rgb <= "100110";
		when "001011100111111" => rgb <= "100110";
		when "001011101000000" => rgb <= "100110";
		when "001011101000001" => rgb <= "000000";
		when "001011101000010" => rgb <= "000000";
		when "001011101000011" => rgb <= "000000";
		when "001011101000100" => rgb <= "000000";
		when "001011101000101" => rgb <= "000000";
		when "001011101000110" => rgb <= "000000";
		when "001011101000111" => rgb <= "000000";
		when "001011101001000" => rgb <= "000000";
		when "001011101010011" => rgb <= "000000";
		when "001011101010100" => rgb <= "100110";
		when "001011101010101" => rgb <= "100110";
		when "001011101010110" => rgb <= "100110";
		when "001011101010111" => rgb <= "000000";
		when "001011101011000" => rgb <= "000000";
		when "001011101011001" => rgb <= "000000";
		when "001011101011010" => rgb <= "000000";
		when "001011101011011" => rgb <= "000000";
		when "001011101011100" => rgb <= "000000";
		when "001011101011101" => rgb <= "100110";
		when "001011101011110" => rgb <= "100110";
		when "001011101011111" => rgb <= "100110";
		when "001011101100000" => rgb <= "000000";
		when "001011101100001" => rgb <= "000000";
		when "001011101100010" => rgb <= "000000";
		when "001011101100011" => rgb <= "000000";
		when "001011101100100" => rgb <= "100110";
		when "001011101100101" => rgb <= "100110";
		when "001011101100110" => rgb <= "100110";
		when "001011101100111" => rgb <= "000000";
		when "001011101101000" => rgb <= "000000";
		when "001011101101001" => rgb <= "000000";
		when "001011101101010" => rgb <= "000000";
		when "001011101101011" => rgb <= "100110";
		when "001011101101100" => rgb <= "100110";
		when "001011101101101" => rgb <= "100110";
		when "001011101101110" => rgb <= "000000";
		when "001011101101111" => rgb <= "000000";
		when "001011101110000" => rgb <= "000000";
		when "001011101110001" => rgb <= "000000";
		when "001011101110010" => rgb <= "100110";
		when "001011101110011" => rgb <= "100110";
		when "001011101110100" => rgb <= "100110";
		when "001011101110101" => rgb <= "000000";
		when "001011101110110" => rgb <= "000000";
		when "001011101110111" => rgb <= "000000";
		when "001011101111000" => rgb <= "000000";
		when "001011101111001" => rgb <= "000000";
		when "001011101111010" => rgb <= "000000";
		when "001011101111011" => rgb <= "000000";
		when "001011101111100" => rgb <= "000000";
		when "001011101111110" => rgb <= "000000";
		when "001011101111111" => rgb <= "100110";
		when "001011110000000" => rgb <= "100110";
		when "001011110000001" => rgb <= "100110";
		when "001011110000010" => rgb <= "100110";
		when "001011110000011" => rgb <= "100110";
		when "001011110000100" => rgb <= "100110";
		when "001011110000101" => rgb <= "100110";
		when "001011110000110" => rgb <= "100110";
		when "001011110000111" => rgb <= "000000";
		when "001011110001000" => rgb <= "000000";
		when "001011110001001" => rgb <= "000000";
		when "001011110001010" => rgb <= "000000";
		when "001100000010010" => rgb <= "000000";
		when "001100000010011" => rgb <= "100110";
		when "001100000010100" => rgb <= "100110";
		when "001100000010101" => rgb <= "100110";
		when "001100000010110" => rgb <= "000000";
		when "001100000010111" => rgb <= "000000";
		when "001100000011000" => rgb <= "000000";
		when "001100000011001" => rgb <= "000000";
		when "001100000011010" => rgb <= "000000";
		when "001100000011011" => rgb <= "000000";
		when "001100000011100" => rgb <= "100110";
		when "001100000011101" => rgb <= "100110";
		when "001100000011110" => rgb <= "100110";
		when "001100000011111" => rgb <= "000000";
		when "001100000100000" => rgb <= "000000";
		when "001100000100001" => rgb <= "100110";
		when "001100000100010" => rgb <= "100110";
		when "001100000100011" => rgb <= "100110";
		when "001100000100100" => rgb <= "000000";
		when "001100000100101" => rgb <= "000000";
		when "001100000100110" => rgb <= "000000";
		when "001100000100111" => rgb <= "000000";
		when "001100000101000" => rgb <= "000000";
		when "001100000101001" => rgb <= "000000";
		when "001100000101010" => rgb <= "100110";
		when "001100000101011" => rgb <= "100110";
		when "001100000101100" => rgb <= "100110";
		when "001100000101101" => rgb <= "000000";
		when "001100000101110" => rgb <= "000000";
		when "001100000101111" => rgb <= "100110";
		when "001100000110000" => rgb <= "100110";
		when "001100000110001" => rgb <= "100110";
		when "001100000110010" => rgb <= "000000";
		when "001100000110011" => rgb <= "000000";
		when "001100000110100" => rgb <= "100110";
		when "001100000110101" => rgb <= "100110";
		when "001100000110110" => rgb <= "100110";
		when "001100000110111" => rgb <= "000000";
		when "001100000111000" => rgb <= "000000";
		when "001100000111001" => rgb <= "100110";
		when "001100000111010" => rgb <= "100110";
		when "001100000111011" => rgb <= "100110";
		when "001100000111100" => rgb <= "000000";
		when "001100000111101" => rgb <= "000000";
		when "001100000111110" => rgb <= "100110";
		when "001100000111111" => rgb <= "100110";
		when "001100001000000" => rgb <= "100110";
		when "001100001000001" => rgb <= "000000";
		when "001100001000010" => rgb <= "000000";
		when "001100001000011" => rgb <= "000000";
		when "001100001000100" => rgb <= "000000";
		when "001100001000101" => rgb <= "000000";
		when "001100001000110" => rgb <= "000000";
		when "001100001000111" => rgb <= "000000";
		when "001100001001000" => rgb <= "000000";
		when "001100001010011" => rgb <= "000000";
		when "001100001010100" => rgb <= "100110";
		when "001100001010101" => rgb <= "100110";
		when "001100001010110" => rgb <= "100110";
		when "001100001010111" => rgb <= "000000";
		when "001100001011000" => rgb <= "000000";
		when "001100001011001" => rgb <= "000000";
		when "001100001011010" => rgb <= "000000";
		when "001100001011011" => rgb <= "000000";
		when "001100001011100" => rgb <= "000000";
		when "001100001011101" => rgb <= "100110";
		when "001100001011110" => rgb <= "100110";
		when "001100001011111" => rgb <= "100110";
		when "001100001100000" => rgb <= "000000";
		when "001100001100001" => rgb <= "000000";
		when "001100001100010" => rgb <= "000000";
		when "001100001100011" => rgb <= "000000";
		when "001100001100100" => rgb <= "100110";
		when "001100001100101" => rgb <= "100110";
		when "001100001100110" => rgb <= "100110";
		when "001100001100111" => rgb <= "000000";
		when "001100001101000" => rgb <= "000000";
		when "001100001101001" => rgb <= "000000";
		when "001100001101010" => rgb <= "000000";
		when "001100001101011" => rgb <= "100110";
		when "001100001101100" => rgb <= "100110";
		when "001100001101101" => rgb <= "100110";
		when "001100001101110" => rgb <= "000000";
		when "001100001101111" => rgb <= "000000";
		when "001100001110000" => rgb <= "000000";
		when "001100001110001" => rgb <= "000000";
		when "001100001110010" => rgb <= "100110";
		when "001100001110011" => rgb <= "100110";
		when "001100001110100" => rgb <= "100110";
		when "001100001110101" => rgb <= "000000";
		when "001100001110110" => rgb <= "000000";
		when "001100001110111" => rgb <= "000000";
		when "001100001111000" => rgb <= "000000";
		when "001100001111001" => rgb <= "000000";
		when "001100001111010" => rgb <= "000000";
		when "001100001111011" => rgb <= "000000";
		when "001100001111100" => rgb <= "000000";
		when "001100001111110" => rgb <= "000000";
		when "001100001111111" => rgb <= "100110";
		when "001100010000000" => rgb <= "100110";
		when "001100010000001" => rgb <= "100110";
		when "001100010000010" => rgb <= "000000";
		when "001100010000011" => rgb <= "000000";
		when "001100010000100" => rgb <= "100110";
		when "001100010000101" => rgb <= "100110";
		when "001100010000110" => rgb <= "100110";
		when "001100010000111" => rgb <= "100110";
		when "001100010001000" => rgb <= "000000";
		when "001100010001001" => rgb <= "000000";
		when "001100010001010" => rgb <= "000000";
		when "001100010001011" => rgb <= "000000";
		when "001100100010010" => rgb <= "000000";
		when "001100100010011" => rgb <= "100110";
		when "001100100010100" => rgb <= "100110";
		when "001100100010101" => rgb <= "100110";
		when "001100100010110" => rgb <= "100110";
		when "001100100010111" => rgb <= "000000";
		when "001100100011000" => rgb <= "000000";
		when "001100100011001" => rgb <= "000000";
		when "001100100011010" => rgb <= "000000";
		when "001100100011011" => rgb <= "000000";
		when "001100100011100" => rgb <= "100110";
		when "001100100011101" => rgb <= "100110";
		when "001100100011110" => rgb <= "100110";
		when "001100100011111" => rgb <= "000000";
		when "001100100100000" => rgb <= "000000";
		when "001100100100001" => rgb <= "100110";
		when "001100100100010" => rgb <= "100110";
		when "001100100100011" => rgb <= "100110";
		when "001100100100100" => rgb <= "000000";
		when "001100100100101" => rgb <= "000000";
		when "001100100100110" => rgb <= "000000";
		when "001100100100111" => rgb <= "000000";
		when "001100100101000" => rgb <= "000000";
		when "001100100101001" => rgb <= "000000";
		when "001100100101010" => rgb <= "100110";
		when "001100100101011" => rgb <= "100110";
		when "001100100101100" => rgb <= "100110";
		when "001100100101101" => rgb <= "000000";
		when "001100100101110" => rgb <= "000000";
		when "001100100101111" => rgb <= "100110";
		when "001100100110000" => rgb <= "100110";
		when "001100100110001" => rgb <= "100110";
		when "001100100110010" => rgb <= "000000";
		when "001100100110011" => rgb <= "000000";
		when "001100100110100" => rgb <= "100110";
		when "001100100110101" => rgb <= "100110";
		when "001100100110110" => rgb <= "100110";
		when "001100100110111" => rgb <= "000000";
		when "001100100111000" => rgb <= "000000";
		when "001100100111001" => rgb <= "100110";
		when "001100100111010" => rgb <= "100110";
		when "001100100111011" => rgb <= "100110";
		when "001100100111100" => rgb <= "000000";
		when "001100100111101" => rgb <= "000000";
		when "001100100111110" => rgb <= "100110";
		when "001100100111111" => rgb <= "100110";
		when "001100101000000" => rgb <= "100110";
		when "001100101000001" => rgb <= "000000";
		when "001100101000010" => rgb <= "000000";
		when "001100101000011" => rgb <= "000000";
		when "001100101000100" => rgb <= "000000";
		when "001100101000101" => rgb <= "000000";
		when "001100101000110" => rgb <= "000000";
		when "001100101000111" => rgb <= "000000";
		when "001100101001000" => rgb <= "000000";
		when "001100101010011" => rgb <= "000000";
		when "001100101010100" => rgb <= "100110";
		when "001100101010101" => rgb <= "100110";
		when "001100101010110" => rgb <= "100110";
		when "001100101010111" => rgb <= "100110";
		when "001100101011000" => rgb <= "000000";
		when "001100101011001" => rgb <= "000000";
		when "001100101011010" => rgb <= "000000";
		when "001100101011011" => rgb <= "000000";
		when "001100101011100" => rgb <= "100110";
		when "001100101011101" => rgb <= "100110";
		when "001100101011110" => rgb <= "100110";
		when "001100101011111" => rgb <= "100110";
		when "001100101100000" => rgb <= "000000";
		when "001100101100001" => rgb <= "000000";
		when "001100101100011" => rgb <= "000000";
		when "001100101100100" => rgb <= "000000";
		when "001100101100101" => rgb <= "100110";
		when "001100101100110" => rgb <= "100110";
		when "001100101100111" => rgb <= "100110";
		when "001100101101000" => rgb <= "100110";
		when "001100101101001" => rgb <= "100110";
		when "001100101101010" => rgb <= "100110";
		when "001100101101011" => rgb <= "100110";
		when "001100101101100" => rgb <= "100110";
		when "001100101101101" => rgb <= "000000";
		when "001100101101110" => rgb <= "000000";
		when "001100101101111" => rgb <= "000000";
		when "001100101110000" => rgb <= "000000";
		when "001100101110001" => rgb <= "000000";
		when "001100101110010" => rgb <= "100110";
		when "001100101110011" => rgb <= "100110";
		when "001100101110100" => rgb <= "100110";
		when "001100101110101" => rgb <= "000000";
		when "001100101110110" => rgb <= "000000";
		when "001100101110111" => rgb <= "000000";
		when "001100101111000" => rgb <= "000000";
		when "001100101111001" => rgb <= "000000";
		when "001100101111010" => rgb <= "000000";
		when "001100101111011" => rgb <= "000000";
		when "001100101111100" => rgb <= "000000";
		when "001100101111110" => rgb <= "000000";
		when "001100101111111" => rgb <= "100110";
		when "001100110000000" => rgb <= "100110";
		when "001100110000001" => rgb <= "100110";
		when "001100110000010" => rgb <= "000000";
		when "001100110000011" => rgb <= "000000";
		when "001100110000100" => rgb <= "000000";
		when "001100110000101" => rgb <= "100110";
		when "001100110000110" => rgb <= "100110";
		when "001100110000111" => rgb <= "100110";
		when "001100110001000" => rgb <= "100110";
		when "001100110001001" => rgb <= "000000";
		when "001100110001010" => rgb <= "000000";
		when "001100110001011" => rgb <= "000000";
		when "001101000010010" => rgb <= "000000";
		when "001101000010011" => rgb <= "100110";
		when "001101000010100" => rgb <= "100110";
		when "001101000010101" => rgb <= "100110";
		when "001101000010110" => rgb <= "100110";
		when "001101000010111" => rgb <= "100110";
		when "001101000011000" => rgb <= "100110";
		when "001101000011001" => rgb <= "100110";
		when "001101000011010" => rgb <= "100110";
		when "001101000011011" => rgb <= "100110";
		when "001101000011100" => rgb <= "100110";
		when "001101000011101" => rgb <= "100110";
		when "001101000011110" => rgb <= "100110";
		when "001101000011111" => rgb <= "000000";
		when "001101000100000" => rgb <= "000000";
		when "001101000100001" => rgb <= "100110";
		when "001101000100010" => rgb <= "100110";
		when "001101000100011" => rgb <= "100110";
		when "001101000100100" => rgb <= "000000";
		when "001101000100101" => rgb <= "000000";
		when "001101000100110" => rgb <= "000000";
		when "001101000100111" => rgb <= "000000";
		when "001101000101000" => rgb <= "000000";
		when "001101000101001" => rgb <= "000000";
		when "001101000101010" => rgb <= "100110";
		when "001101000101011" => rgb <= "100110";
		when "001101000101100" => rgb <= "100110";
		when "001101000101101" => rgb <= "000000";
		when "001101000101110" => rgb <= "000000";
		when "001101000101111" => rgb <= "100110";
		when "001101000110000" => rgb <= "100110";
		when "001101000110001" => rgb <= "100110";
		when "001101000110010" => rgb <= "000000";
		when "001101000110011" => rgb <= "000000";
		when "001101000110100" => rgb <= "000000";
		when "001101000110101" => rgb <= "000000";
		when "001101000110110" => rgb <= "000000";
		when "001101000110111" => rgb <= "000000";
		when "001101000111000" => rgb <= "000000";
		when "001101000111001" => rgb <= "100110";
		when "001101000111010" => rgb <= "100110";
		when "001101000111011" => rgb <= "100110";
		when "001101000111100" => rgb <= "000000";
		when "001101000111101" => rgb <= "000000";
		when "001101000111110" => rgb <= "100110";
		when "001101000111111" => rgb <= "100110";
		when "001101001000000" => rgb <= "100110";
		when "001101001000001" => rgb <= "100110";
		when "001101001000010" => rgb <= "100110";
		when "001101001000011" => rgb <= "100110";
		when "001101001000100" => rgb <= "100110";
		when "001101001000101" => rgb <= "100110";
		when "001101001000110" => rgb <= "100110";
		when "001101001000111" => rgb <= "100110";
		when "001101001001000" => rgb <= "000000";
		when "001101001001001" => rgb <= "000000";
		when "001101001001010" => rgb <= "000000";
		when "001101001010011" => rgb <= "000000";
		when "001101001010100" => rgb <= "000000";
		when "001101001010101" => rgb <= "100110";
		when "001101001010110" => rgb <= "100110";
		when "001101001010111" => rgb <= "100110";
		when "001101001011000" => rgb <= "100110";
		when "001101001011001" => rgb <= "100110";
		when "001101001011010" => rgb <= "100110";
		when "001101001011011" => rgb <= "100110";
		when "001101001011100" => rgb <= "100110";
		when "001101001011101" => rgb <= "100110";
		when "001101001011110" => rgb <= "100110";
		when "001101001011111" => rgb <= "000000";
		when "001101001100000" => rgb <= "000000";
		when "001101001100001" => rgb <= "000000";
		when "001101001100011" => rgb <= "000000";
		when "001101001100100" => rgb <= "000000";
		when "001101001100101" => rgb <= "100110";
		when "001101001100110" => rgb <= "100110";
		when "001101001100111" => rgb <= "100110";
		when "001101001101000" => rgb <= "100110";
		when "001101001101001" => rgb <= "100110";
		when "001101001101010" => rgb <= "100110";
		when "001101001101011" => rgb <= "100110";
		when "001101001101100" => rgb <= "100110";
		when "001101001101101" => rgb <= "000000";
		when "001101001101110" => rgb <= "000000";
		when "001101001101111" => rgb <= "000000";
		when "001101001110001" => rgb <= "000000";
		when "001101001110010" => rgb <= "100110";
		when "001101001110011" => rgb <= "100110";
		when "001101001110100" => rgb <= "100110";
		when "001101001110101" => rgb <= "100110";
		when "001101001110110" => rgb <= "100110";
		when "001101001110111" => rgb <= "100110";
		when "001101001111000" => rgb <= "100110";
		when "001101001111001" => rgb <= "100110";
		when "001101001111010" => rgb <= "100110";
		when "001101001111011" => rgb <= "100110";
		when "001101001111100" => rgb <= "000000";
		when "001101001111101" => rgb <= "000000";
		when "001101001111110" => rgb <= "000000";
		when "001101001111111" => rgb <= "100110";
		when "001101010000000" => rgb <= "100110";
		when "001101010000001" => rgb <= "100110";
		when "001101010000010" => rgb <= "000000";
		when "001101010000011" => rgb <= "000000";
		when "001101010000100" => rgb <= "000000";
		when "001101010000101" => rgb <= "000000";
		when "001101010000110" => rgb <= "100110";
		when "001101010000111" => rgb <= "100110";
		when "001101010001000" => rgb <= "100110";
		when "001101010001001" => rgb <= "000000";
		when "001101010001010" => rgb <= "000000";
		when "001101010001011" => rgb <= "000000";
		when "001101100010010" => rgb <= "000000";
		when "001101100010011" => rgb <= "000000";
		when "001101100010100" => rgb <= "100110";
		when "001101100010101" => rgb <= "100110";
		when "001101100010110" => rgb <= "100110";
		when "001101100010111" => rgb <= "100110";
		when "001101100011000" => rgb <= "100110";
		when "001101100011001" => rgb <= "100110";
		when "001101100011010" => rgb <= "100110";
		when "001101100011011" => rgb <= "100110";
		when "001101100011100" => rgb <= "100110";
		when "001101100011101" => rgb <= "100110";
		when "001101100011110" => rgb <= "100110";
		when "001101100011111" => rgb <= "000000";
		when "001101100100000" => rgb <= "000000";
		when "001101100100001" => rgb <= "100110";
		when "001101100100010" => rgb <= "100110";
		when "001101100100011" => rgb <= "100110";
		when "001101100100100" => rgb <= "000000";
		when "001101100100101" => rgb <= "000000";
		when "001101100100110" => rgb <= "000000";
		when "001101100101001" => rgb <= "000000";
		when "001101100101010" => rgb <= "100110";
		when "001101100101011" => rgb <= "100110";
		when "001101100101100" => rgb <= "100110";
		when "001101100101101" => rgb <= "000000";
		when "001101100101110" => rgb <= "000000";
		when "001101100101111" => rgb <= "100110";
		when "001101100110000" => rgb <= "100110";
		when "001101100110001" => rgb <= "100110";
		when "001101100110010" => rgb <= "000000";
		when "001101100110011" => rgb <= "000000";
		when "001101100110100" => rgb <= "000000";
		when "001101100110101" => rgb <= "000000";
		when "001101100110110" => rgb <= "000000";
		when "001101100110111" => rgb <= "000000";
		when "001101100111000" => rgb <= "000000";
		when "001101100111001" => rgb <= "100110";
		when "001101100111010" => rgb <= "100110";
		when "001101100111011" => rgb <= "100110";
		when "001101100111100" => rgb <= "000000";
		when "001101100111101" => rgb <= "000000";
		when "001101100111110" => rgb <= "100110";
		when "001101100111111" => rgb <= "100110";
		when "001101101000000" => rgb <= "100110";
		when "001101101000001" => rgb <= "100110";
		when "001101101000010" => rgb <= "100110";
		when "001101101000011" => rgb <= "100110";
		when "001101101000100" => rgb <= "100110";
		when "001101101000101" => rgb <= "100110";
		when "001101101000110" => rgb <= "100110";
		when "001101101000111" => rgb <= "100110";
		when "001101101001000" => rgb <= "000000";
		when "001101101001001" => rgb <= "000000";
		when "001101101001010" => rgb <= "000000";
		when "001101101010011" => rgb <= "000000";
		when "001101101010100" => rgb <= "000000";
		when "001101101010101" => rgb <= "100110";
		when "001101101010110" => rgb <= "100110";
		when "001101101010111" => rgb <= "100110";
		when "001101101011000" => rgb <= "100110";
		when "001101101011001" => rgb <= "100110";
		when "001101101011010" => rgb <= "100110";
		when "001101101011011" => rgb <= "100110";
		when "001101101011100" => rgb <= "100110";
		when "001101101011101" => rgb <= "100110";
		when "001101101011110" => rgb <= "100110";
		when "001101101011111" => rgb <= "000000";
		when "001101101100000" => rgb <= "000000";
		when "001101101100001" => rgb <= "000000";
		when "001101101100100" => rgb <= "000000";
		when "001101101100101" => rgb <= "000000";
		when "001101101100110" => rgb <= "000000";
		when "001101101100111" => rgb <= "100110";
		when "001101101101000" => rgb <= "100110";
		when "001101101101001" => rgb <= "100110";
		when "001101101101010" => rgb <= "100110";
		when "001101101101011" => rgb <= "000000";
		when "001101101101100" => rgb <= "000000";
		when "001101101101101" => rgb <= "000000";
		when "001101101101110" => rgb <= "000000";
		when "001101101110001" => rgb <= "000000";
		when "001101101110010" => rgb <= "100110";
		when "001101101110011" => rgb <= "100110";
		when "001101101110100" => rgb <= "100110";
		when "001101101110101" => rgb <= "100110";
		when "001101101110110" => rgb <= "100110";
		when "001101101110111" => rgb <= "100110";
		when "001101101111000" => rgb <= "100110";
		when "001101101111001" => rgb <= "100110";
		when "001101101111010" => rgb <= "100110";
		when "001101101111011" => rgb <= "100110";
		when "001101101111100" => rgb <= "000000";
		when "001101101111101" => rgb <= "000000";
		when "001101101111110" => rgb <= "000000";
		when "001101101111111" => rgb <= "100110";
		when "001101110000000" => rgb <= "100110";
		when "001101110000001" => rgb <= "100110";
		when "001101110000010" => rgb <= "000000";
		when "001101110000011" => rgb <= "000000";
		when "001101110000100" => rgb <= "000000";
		when "001101110000101" => rgb <= "000000";
		when "001101110000110" => rgb <= "100110";
		when "001101110000111" => rgb <= "100110";
		when "001101110001000" => rgb <= "100110";
		when "001101110001001" => rgb <= "000000";
		when "001101110001010" => rgb <= "000000";
		when "001101110001011" => rgb <= "000000";
		when "001110000010011" => rgb <= "000000";
		when "001110000010100" => rgb <= "000000";
		when "001110000010101" => rgb <= "000000";
		when "001110000010110" => rgb <= "100110";
		when "001110000010111" => rgb <= "100110";
		when "001110000011000" => rgb <= "100110";
		when "001110000011001" => rgb <= "100110";
		when "001110000011010" => rgb <= "100110";
		when "001110000011011" => rgb <= "100110";
		when "001110000011100" => rgb <= "100110";
		when "001110000011101" => rgb <= "100110";
		when "001110000011110" => rgb <= "100110";
		when "001110000011111" => rgb <= "000000";
		when "001110000100000" => rgb <= "000000";
		when "001110000100001" => rgb <= "100110";
		when "001110000100010" => rgb <= "100110";
		when "001110000100011" => rgb <= "100110";
		when "001110000100100" => rgb <= "000000";
		when "001110000100101" => rgb <= "000000";
		when "001110000100110" => rgb <= "000000";
		when "001110000101001" => rgb <= "000000";
		when "001110000101010" => rgb <= "100110";
		when "001110000101011" => rgb <= "100110";
		when "001110000101100" => rgb <= "100110";
		when "001110000101101" => rgb <= "000000";
		when "001110000101110" => rgb <= "000000";
		when "001110000101111" => rgb <= "100110";
		when "001110000110000" => rgb <= "100110";
		when "001110000110001" => rgb <= "100110";
		when "001110000110010" => rgb <= "000000";
		when "001110000110011" => rgb <= "000000";
		when "001110000110101" => rgb <= "000000";
		when "001110000110110" => rgb <= "000000";
		when "001110000110111" => rgb <= "000000";
		when "001110000111000" => rgb <= "000000";
		when "001110000111001" => rgb <= "100110";
		when "001110000111010" => rgb <= "100110";
		when "001110000111011" => rgb <= "100110";
		when "001110000111100" => rgb <= "000000";
		when "001110000111101" => rgb <= "000000";
		when "001110000111110" => rgb <= "100110";
		when "001110000111111" => rgb <= "100110";
		when "001110001000000" => rgb <= "100110";
		when "001110001000001" => rgb <= "100110";
		when "001110001000010" => rgb <= "100110";
		when "001110001000011" => rgb <= "100110";
		when "001110001000100" => rgb <= "100110";
		when "001110001000101" => rgb <= "100110";
		when "001110001000110" => rgb <= "100110";
		when "001110001000111" => rgb <= "100110";
		when "001110001001000" => rgb <= "000000";
		when "001110001001001" => rgb <= "000000";
		when "001110001001010" => rgb <= "000000";
		when "001110001010011" => rgb <= "000000";
		when "001110001010100" => rgb <= "000000";
		when "001110001010101" => rgb <= "000000";
		when "001110001010110" => rgb <= "000000";
		when "001110001010111" => rgb <= "100110";
		when "001110001011000" => rgb <= "100110";
		when "001110001011001" => rgb <= "100110";
		when "001110001011010" => rgb <= "100110";
		when "001110001011011" => rgb <= "100110";
		when "001110001011100" => rgb <= "100110";
		when "001110001011101" => rgb <= "000000";
		when "001110001011110" => rgb <= "000000";
		when "001110001011111" => rgb <= "000000";
		when "001110001100000" => rgb <= "000000";
		when "001110001100001" => rgb <= "000000";
		when "001110001100101" => rgb <= "000000";
		when "001110001100110" => rgb <= "000000";
		when "001110001100111" => rgb <= "000000";
		when "001110001101000" => rgb <= "100110";
		when "001110001101001" => rgb <= "100110";
		when "001110001101010" => rgb <= "000000";
		when "001110001101011" => rgb <= "000000";
		when "001110001101100" => rgb <= "000000";
		when "001110001101101" => rgb <= "000000";
		when "001110001110001" => rgb <= "000000";
		when "001110001110010" => rgb <= "100110";
		when "001110001110011" => rgb <= "100110";
		when "001110001110100" => rgb <= "100110";
		when "001110001110101" => rgb <= "100110";
		when "001110001110110" => rgb <= "100110";
		when "001110001110111" => rgb <= "100110";
		when "001110001111000" => rgb <= "100110";
		when "001110001111001" => rgb <= "100110";
		when "001110001111010" => rgb <= "100110";
		when "001110001111011" => rgb <= "100110";
		when "001110001111100" => rgb <= "000000";
		when "001110001111101" => rgb <= "000000";
		when "001110001111110" => rgb <= "000000";
		when "001110001111111" => rgb <= "100110";
		when "001110010000000" => rgb <= "100110";
		when "001110010000001" => rgb <= "100110";
		when "001110010000010" => rgb <= "000000";
		when "001110010000011" => rgb <= "000000";
		when "001110010000100" => rgb <= "000000";
		when "001110010000101" => rgb <= "000000";
		when "001110010000110" => rgb <= "100110";
		when "001110010000111" => rgb <= "100110";
		when "001110010001000" => rgb <= "100110";
		when "001110010001001" => rgb <= "000000";
		when "001110010001010" => rgb <= "000000";
		when "001110010001011" => rgb <= "000000";
		when "001110100010100" => rgb <= "000000";
		when "001110100010101" => rgb <= "000000";
		when "001110100010110" => rgb <= "000000";
		when "001110100010111" => rgb <= "000000";
		when "001110100011000" => rgb <= "000000";
		when "001110100011001" => rgb <= "000000";
		when "001110100011010" => rgb <= "000000";
		when "001110100011011" => rgb <= "000000";
		when "001110100011100" => rgb <= "000000";
		when "001110100011101" => rgb <= "000000";
		when "001110100011110" => rgb <= "000000";
		when "001110100011111" => rgb <= "000000";
		when "001110100100000" => rgb <= "000000";
		when "001110100100001" => rgb <= "000000";
		when "001110100100010" => rgb <= "000000";
		when "001110100100011" => rgb <= "000000";
		when "001110100100100" => rgb <= "000000";
		when "001110100100101" => rgb <= "000000";
		when "001110100100110" => rgb <= "000000";
		when "001110100101001" => rgb <= "000000";
		when "001110100101010" => rgb <= "000000";
		when "001110100101011" => rgb <= "000000";
		when "001110100101100" => rgb <= "000000";
		when "001110100101101" => rgb <= "000000";
		when "001110100101110" => rgb <= "000000";
		when "001110100101111" => rgb <= "000000";
		when "001110100110000" => rgb <= "000000";
		when "001110100110001" => rgb <= "000000";
		when "001110100110010" => rgb <= "000000";
		when "001110100110011" => rgb <= "000000";
		when "001110100110110" => rgb <= "000000";
		when "001110100110111" => rgb <= "000000";
		when "001110100111000" => rgb <= "000000";
		when "001110100111001" => rgb <= "000000";
		when "001110100111010" => rgb <= "000000";
		when "001110100111011" => rgb <= "000000";
		when "001110100111100" => rgb <= "000000";
		when "001110100111101" => rgb <= "000000";
		when "001110100111110" => rgb <= "000000";
		when "001110100111111" => rgb <= "000000";
		when "001110101000000" => rgb <= "000000";
		when "001110101000001" => rgb <= "000000";
		when "001110101000010" => rgb <= "000000";
		when "001110101000011" => rgb <= "000000";
		when "001110101000100" => rgb <= "000000";
		when "001110101000101" => rgb <= "000000";
		when "001110101000110" => rgb <= "000000";
		when "001110101000111" => rgb <= "000000";
		when "001110101001000" => rgb <= "000000";
		when "001110101001001" => rgb <= "000000";
		when "001110101001010" => rgb <= "000000";
		when "001110101010100" => rgb <= "000000";
		when "001110101010101" => rgb <= "000000";
		when "001110101010110" => rgb <= "000000";
		when "001110101010111" => rgb <= "000000";
		when "001110101011000" => rgb <= "000000";
		when "001110101011001" => rgb <= "000000";
		when "001110101011010" => rgb <= "000000";
		when "001110101011011" => rgb <= "000000";
		when "001110101011100" => rgb <= "000000";
		when "001110101011101" => rgb <= "000000";
		when "001110101011110" => rgb <= "000000";
		when "001110101011111" => rgb <= "000000";
		when "001110101100000" => rgb <= "000000";
		when "001110101100101" => rgb <= "000000";
		when "001110101100110" => rgb <= "000000";
		when "001110101100111" => rgb <= "000000";
		when "001110101101000" => rgb <= "000000";
		when "001110101101001" => rgb <= "000000";
		when "001110101101010" => rgb <= "000000";
		when "001110101101011" => rgb <= "000000";
		when "001110101101100" => rgb <= "000000";
		when "001110101110001" => rgb <= "000000";
		when "001110101110010" => rgb <= "000000";
		when "001110101110011" => rgb <= "000000";
		when "001110101110100" => rgb <= "000000";
		when "001110101110101" => rgb <= "000000";
		when "001110101110110" => rgb <= "000000";
		when "001110101110111" => rgb <= "000000";
		when "001110101111000" => rgb <= "000000";
		when "001110101111001" => rgb <= "000000";
		when "001110101111010" => rgb <= "000000";
		when "001110101111011" => rgb <= "000000";
		when "001110101111100" => rgb <= "000000";
		when "001110101111101" => rgb <= "000000";
		when "001110101111110" => rgb <= "000000";
		when "001110101111111" => rgb <= "000000";
		when "001110110000000" => rgb <= "000000";
		when "001110110000001" => rgb <= "000000";
		when "001110110000010" => rgb <= "000000";
		when "001110110000011" => rgb <= "000000";
		when "001110110000101" => rgb <= "000000";
		when "001110110000110" => rgb <= "000000";
		when "001110110000111" => rgb <= "000000";
		when "001110110001000" => rgb <= "000000";
		when "001110110001001" => rgb <= "000000";
		when "001110110001010" => rgb <= "000000";
		when "001110110001011" => rgb <= "000000";
		when "001111000010100" => rgb <= "000000";
		when "001111000010101" => rgb <= "000000";
		when "001111000010110" => rgb <= "000000";
		when "001111000010111" => rgb <= "000000";
		when "001111000011000" => rgb <= "000000";
		when "001111000011001" => rgb <= "000000";
		when "001111000011010" => rgb <= "000000";
		when "001111000011011" => rgb <= "000000";
		when "001111000011100" => rgb <= "000000";
		when "001111000011101" => rgb <= "000000";
		when "001111000011110" => rgb <= "000000";
		when "001111000011111" => rgb <= "000000";
		when "001111000100000" => rgb <= "000000";
		when "001111000100010" => rgb <= "000000";
		when "001111000100011" => rgb <= "000000";
		when "001111000100100" => rgb <= "000000";
		when "001111000100101" => rgb <= "000000";
		when "001111000100110" => rgb <= "000000";
		when "001111000101010" => rgb <= "000000";
		when "001111000101011" => rgb <= "000000";
		when "001111000101100" => rgb <= "000000";
		when "001111000101101" => rgb <= "000000";
		when "001111000101110" => rgb <= "000000";
		when "001111000110000" => rgb <= "000000";
		when "001111000110001" => rgb <= "000000";
		when "001111000110010" => rgb <= "000000";
		when "001111000110011" => rgb <= "000000";
		when "001111000111001" => rgb <= "000000";
		when "001111000111010" => rgb <= "000000";
		when "001111000111011" => rgb <= "000000";
		when "001111000111100" => rgb <= "000000";
		when "001111000111101" => rgb <= "000000";
		when "001111000111111" => rgb <= "000000";
		when "001111001000000" => rgb <= "000000";
		when "001111001000001" => rgb <= "000000";
		when "001111001000010" => rgb <= "000000";
		when "001111001000011" => rgb <= "000000";
		when "001111001000100" => rgb <= "000000";
		when "001111001000101" => rgb <= "000000";
		when "001111001000110" => rgb <= "000000";
		when "001111001000111" => rgb <= "000000";
		when "001111001001000" => rgb <= "000000";
		when "001111001001001" => rgb <= "000000";
		when "001111001001010" => rgb <= "000000";
		when "001111001010100" => rgb <= "000000";
		when "001111001010101" => rgb <= "000000";
		when "001111001010110" => rgb <= "000000";
		when "001111001010111" => rgb <= "000000";
		when "001111001011000" => rgb <= "000000";
		when "001111001011001" => rgb <= "000000";
		when "001111001011010" => rgb <= "000000";
		when "001111001011011" => rgb <= "000000";
		when "001111001011100" => rgb <= "000000";
		when "001111001011101" => rgb <= "000000";
		when "001111001011110" => rgb <= "000000";
		when "001111001011111" => rgb <= "000000";
		when "001111001100111" => rgb <= "000000";
		when "001111001101000" => rgb <= "000000";
		when "001111001101001" => rgb <= "000000";
		when "001111001101010" => rgb <= "000000";
		when "001111001110011" => rgb <= "000000";
		when "001111001110100" => rgb <= "000000";
		when "001111001110101" => rgb <= "000000";
		when "001111001110110" => rgb <= "000000";
		when "001111001110111" => rgb <= "000000";
		when "001111001111000" => rgb <= "000000";
		when "001111001111001" => rgb <= "000000";
		when "001111001111010" => rgb <= "000000";
		when "001111001111011" => rgb <= "000000";
		when "001111001111100" => rgb <= "000000";
		when "001111001111101" => rgb <= "000000";
		when "001111001111110" => rgb <= "000000";
		when "001111010000000" => rgb <= "000000";
		when "001111010000001" => rgb <= "000000";
		when "001111010000010" => rgb <= "000000";
		when "001111010000011" => rgb <= "000000";
		when "001111010000111" => rgb <= "000000";
		when "001111010001000" => rgb <= "000000";
		when "001111010001001" => rgb <= "000000";
		when "001111010001010" => rgb <= "000000";
		when "001111010001011" => rgb <= "000000";
		when "001111100010101" => rgb <= "000000";
		when "001111100010110" => rgb <= "000000";
		when "001111100010111" => rgb <= "000000";
		when "001111100011000" => rgb <= "000000";
		when "001111100011001" => rgb <= "000000";
		when "001111100011010" => rgb <= "000000";
		when "001111100011011" => rgb <= "000000";
		when "001111100011100" => rgb <= "000000";
		when "001111100011101" => rgb <= "000000";
		when "001111100011110" => rgb <= "000000";
		when "001111100011111" => rgb <= "000000";
		when "001111100100000" => rgb <= "000000";
		when "001111100100010" => rgb <= "000000";
		when "001111100100011" => rgb <= "000000";
		when "001111100100100" => rgb <= "000000";
		when "001111100100101" => rgb <= "000000";
		when "001111100100110" => rgb <= "000000";
		when "001111100101010" => rgb <= "000000";
		when "001111100101011" => rgb <= "000000";
		when "001111100101100" => rgb <= "000000";
		when "001111100101101" => rgb <= "000000";
		when "001111100101110" => rgb <= "000000";
		when "001111100110000" => rgb <= "000000";
		when "001111100110001" => rgb <= "000000";
		when "001111100110010" => rgb <= "000000";
		when "001111100110011" => rgb <= "000000";
		when "001111100111001" => rgb <= "000000";
		when "001111100111010" => rgb <= "000000";
		when "001111100111011" => rgb <= "000000";
		when "001111100111100" => rgb <= "000000";
		when "001111100111101" => rgb <= "000000";
		when "001111100111111" => rgb <= "000000";
		when "001111101000000" => rgb <= "000000";
		when "001111101000001" => rgb <= "000000";
		when "001111101000010" => rgb <= "000000";
		when "001111101000011" => rgb <= "000000";
		when "001111101000100" => rgb <= "000000";
		when "001111101000101" => rgb <= "000000";
		when "001111101000110" => rgb <= "000000";
		when "001111101000111" => rgb <= "000000";
		when "001111101001000" => rgb <= "000000";
		when "001111101001001" => rgb <= "000000";
		when "001111101001010" => rgb <= "000000";
		when "001111101010110" => rgb <= "000000";
		when "001111101010111" => rgb <= "000000";
		when "001111101011000" => rgb <= "000000";
		when "001111101011001" => rgb <= "000000";
		when "001111101011010" => rgb <= "000000";
		when "001111101011011" => rgb <= "000000";
		when "001111101011100" => rgb <= "000000";
		when "001111101011101" => rgb <= "000000";
		when "001111101100111" => rgb <= "000000";
		when "001111101101000" => rgb <= "000000";
		when "001111101101001" => rgb <= "000000";
		when "001111101101010" => rgb <= "000000";
		when "001111101110011" => rgb <= "000000";
		when "001111101110100" => rgb <= "000000";
		when "001111101110101" => rgb <= "000000";
		when "001111101110110" => rgb <= "000000";
		when "001111101110111" => rgb <= "000000";
		when "001111101111000" => rgb <= "000000";
		when "001111101111001" => rgb <= "000000";
		when "001111101111010" => rgb <= "000000";
		when "001111101111011" => rgb <= "000000";
		when "001111101111100" => rgb <= "000000";
		when "001111101111101" => rgb <= "000000";
		when "001111101111110" => rgb <= "000000";
		when "001111110000000" => rgb <= "000000";
		when "001111110000001" => rgb <= "000000";
		when "001111110000010" => rgb <= "000000";
		when "001111110000011" => rgb <= "000000";
		when "001111110000111" => rgb <= "000000";
		when "001111110001000" => rgb <= "000000";
		when "001111110001001" => rgb <= "000000";
		when "001111110001010" => rgb <= "000000";
		when "001111110001011" => rgb <= "000000";
		when others => rgb <= "111111"; 
	end case;
end if;
end process;
	addressOut <= address;
end;
